magic
tech scmos
timestamp 1732102314
<< nwell >>
rect 488 221 612 258
rect 253 177 337 214
rect 488 132 612 169
rect 253 94 277 131
rect 631 86 755 123
rect 1225 97 1309 134
rect 0 44 117 71
rect 243 27 305 64
rect 488 49 550 86
rect 1225 14 1249 51
rect 0 -30 117 -3
rect 253 -47 337 -10
rect 488 -42 674 -5
rect 1225 -53 1309 -16
rect 1486 -27 1603 0
rect 0 -104 117 -77
rect 253 -130 277 -93
rect 488 -139 612 -102
rect 718 -126 904 -89
rect 1225 -136 1249 -99
rect 1486 -101 1603 -74
rect 0 -178 117 -151
rect 243 -197 305 -160
rect 488 -224 550 -187
rect 1225 -203 1309 -166
rect 1486 -175 1603 -148
rect 0 -252 117 -225
rect 253 -271 337 -234
rect 1486 -249 1603 -222
rect 1225 -286 1249 -249
rect 0 -326 117 -299
rect 253 -354 277 -317
rect 488 -336 736 -299
rect 1225 -353 1309 -316
rect 1486 -323 1603 -296
rect 0 -400 117 -373
rect 243 -421 305 -384
rect 488 -436 674 -399
rect 1225 -436 1249 -399
rect 0 -474 117 -447
rect 253 -495 337 -458
rect 488 -536 612 -499
rect 796 -518 1044 -481
rect 253 -578 277 -541
rect 243 -645 305 -608
rect 488 -636 550 -599
<< ntransistor >>
rect 499 195 501 205
rect 513 195 515 205
rect 537 195 539 205
rect 561 189 563 199
rect 575 189 577 199
rect 599 189 601 199
rect 264 158 266 168
rect 499 106 501 116
rect 513 106 515 116
rect 537 106 539 116
rect 561 106 563 116
rect 575 106 577 116
rect 599 106 601 116
rect 264 75 266 85
rect 288 75 290 85
rect 305 75 307 85
rect 318 75 320 85
rect 335 75 337 85
rect 1236 78 1238 88
rect 642 54 644 64
rect 656 54 658 64
rect 680 54 682 64
rect 704 54 706 64
rect 718 54 720 64
rect 742 54 744 64
rect 11 10 13 20
rect 42 10 44 20
rect 57 10 59 20
rect 73 10 75 20
rect 88 10 90 20
rect 104 10 106 20
rect 499 23 501 33
rect 513 23 515 33
rect 537 23 539 33
rect 254 1 256 11
rect 268 1 270 11
rect 292 1 294 11
rect 1236 -5 1238 5
rect 1260 -5 1262 5
rect 1277 -5 1279 5
rect 1290 -5 1292 5
rect 1307 -5 1309 5
rect 11 -64 13 -54
rect 42 -64 44 -54
rect 57 -64 59 -54
rect 73 -64 75 -54
rect 88 -64 90 -54
rect 104 -64 106 -54
rect 264 -66 266 -56
rect 11 -138 13 -128
rect 42 -138 44 -128
rect 57 -138 59 -128
rect 73 -138 75 -128
rect 88 -138 90 -128
rect 104 -138 106 -128
rect 499 -68 501 -58
rect 513 -68 515 -58
rect 537 -68 539 -58
rect 561 -68 563 -58
rect 575 -68 577 -58
rect 599 -68 601 -58
rect 623 -68 625 -58
rect 637 -68 639 -58
rect 661 -68 663 -58
rect 1236 -72 1238 -62
rect 264 -149 266 -139
rect 288 -149 290 -139
rect 305 -149 307 -139
rect 318 -149 320 -139
rect 335 -149 337 -139
rect 1497 -61 1499 -51
rect 1528 -61 1530 -51
rect 1543 -61 1545 -51
rect 1559 -61 1561 -51
rect 1574 -61 1576 -51
rect 1590 -61 1592 -51
rect 1497 -135 1499 -125
rect 1528 -135 1530 -125
rect 1543 -135 1545 -125
rect 1559 -135 1561 -125
rect 1574 -135 1576 -125
rect 1590 -135 1592 -125
rect 499 -165 501 -155
rect 513 -165 515 -155
rect 537 -165 539 -155
rect 561 -165 563 -155
rect 575 -165 577 -155
rect 599 -165 601 -155
rect 729 -158 731 -148
rect 743 -158 745 -148
rect 767 -158 769 -148
rect 791 -158 793 -148
rect 805 -158 807 -148
rect 829 -158 831 -148
rect 853 -158 855 -148
rect 867 -158 869 -148
rect 891 -158 893 -148
rect 1236 -155 1238 -145
rect 1260 -155 1262 -145
rect 1277 -155 1279 -145
rect 1290 -155 1292 -145
rect 1307 -155 1309 -145
rect 11 -212 13 -202
rect 42 -212 44 -202
rect 57 -212 59 -202
rect 73 -212 75 -202
rect 88 -212 90 -202
rect 104 -212 106 -202
rect 254 -223 256 -213
rect 268 -223 270 -213
rect 292 -223 294 -213
rect 1236 -222 1238 -212
rect 499 -250 501 -240
rect 513 -250 515 -240
rect 537 -250 539 -240
rect 11 -286 13 -276
rect 42 -286 44 -276
rect 57 -286 59 -276
rect 73 -286 75 -276
rect 88 -286 90 -276
rect 104 -286 106 -276
rect 264 -290 266 -280
rect 11 -360 13 -350
rect 42 -360 44 -350
rect 57 -360 59 -350
rect 73 -360 75 -350
rect 88 -360 90 -350
rect 104 -360 106 -350
rect 1497 -209 1499 -199
rect 1528 -209 1530 -199
rect 1543 -209 1545 -199
rect 1559 -209 1561 -199
rect 1574 -209 1576 -199
rect 1590 -209 1592 -199
rect 1497 -283 1499 -273
rect 1528 -283 1530 -273
rect 1543 -283 1545 -273
rect 1559 -283 1561 -273
rect 1574 -283 1576 -273
rect 1590 -283 1592 -273
rect 1236 -305 1238 -295
rect 1260 -305 1262 -295
rect 1277 -305 1279 -295
rect 1290 -305 1292 -295
rect 1307 -305 1309 -295
rect 499 -362 501 -352
rect 513 -362 515 -352
rect 537 -362 539 -352
rect 561 -362 563 -352
rect 575 -362 577 -352
rect 599 -362 601 -352
rect 623 -362 625 -352
rect 637 -362 639 -352
rect 661 -362 663 -352
rect 685 -362 687 -352
rect 699 -362 701 -352
rect 723 -362 725 -352
rect 264 -373 266 -363
rect 288 -373 290 -363
rect 305 -373 307 -363
rect 318 -373 320 -363
rect 335 -373 337 -363
rect 1236 -372 1238 -362
rect 11 -434 13 -424
rect 42 -434 44 -424
rect 57 -434 59 -424
rect 73 -434 75 -424
rect 88 -434 90 -424
rect 104 -434 106 -424
rect 254 -447 256 -437
rect 268 -447 270 -437
rect 292 -447 294 -437
rect 1497 -357 1499 -347
rect 1528 -357 1530 -347
rect 1543 -357 1545 -347
rect 1559 -357 1561 -347
rect 1574 -357 1576 -347
rect 1590 -357 1592 -347
rect 499 -462 501 -452
rect 513 -462 515 -452
rect 537 -462 539 -452
rect 561 -462 563 -452
rect 575 -462 577 -452
rect 599 -462 601 -452
rect 623 -462 625 -452
rect 637 -462 639 -452
rect 661 -462 663 -452
rect 1236 -455 1238 -445
rect 1260 -455 1262 -445
rect 1277 -455 1279 -445
rect 1290 -455 1292 -445
rect 1307 -455 1309 -445
rect 11 -508 13 -498
rect 42 -508 44 -498
rect 57 -508 59 -498
rect 73 -508 75 -498
rect 88 -508 90 -498
rect 104 -508 106 -498
rect 264 -514 266 -504
rect 807 -550 809 -540
rect 821 -550 823 -540
rect 845 -550 847 -540
rect 869 -550 871 -540
rect 883 -550 885 -540
rect 907 -550 909 -540
rect 931 -550 933 -540
rect 945 -550 947 -540
rect 969 -550 971 -540
rect 993 -550 995 -540
rect 1007 -550 1009 -540
rect 1031 -550 1033 -540
rect 499 -562 501 -552
rect 513 -562 515 -552
rect 537 -562 539 -552
rect 561 -562 563 -552
rect 575 -562 577 -552
rect 599 -562 601 -552
rect 264 -597 266 -587
rect 288 -597 290 -587
rect 305 -597 307 -587
rect 318 -597 320 -587
rect 335 -597 337 -587
rect 254 -671 256 -661
rect 268 -671 270 -661
rect 292 -671 294 -661
rect 499 -662 501 -652
rect 513 -662 515 -652
rect 537 -662 539 -652
<< ptransistor >>
rect 499 227 501 247
rect 513 227 515 247
rect 537 227 539 247
rect 561 227 563 247
rect 575 227 577 247
rect 599 227 601 247
rect 264 183 266 203
rect 288 183 290 203
rect 302 183 304 203
rect 310 183 312 203
rect 324 183 326 203
rect 264 100 266 120
rect 499 138 501 158
rect 513 138 515 158
rect 537 138 539 158
rect 561 138 563 158
rect 575 138 577 158
rect 599 138 601 158
rect 642 92 644 112
rect 656 92 658 112
rect 680 92 682 112
rect 704 92 706 112
rect 718 92 720 112
rect 742 92 744 112
rect 1236 103 1238 123
rect 1260 103 1262 123
rect 1274 103 1276 123
rect 1282 103 1284 123
rect 1296 103 1298 123
rect 11 50 13 60
rect 26 50 28 60
rect 42 50 44 60
rect 73 50 75 60
rect 104 50 106 60
rect 499 55 501 75
rect 513 55 515 75
rect 537 55 539 75
rect 254 33 256 53
rect 268 33 270 53
rect 292 33 294 53
rect 1236 20 1238 40
rect 11 -24 13 -14
rect 26 -24 28 -14
rect 42 -24 44 -14
rect 73 -24 75 -14
rect 104 -24 106 -14
rect 264 -41 266 -21
rect 288 -41 290 -21
rect 302 -41 304 -21
rect 310 -41 312 -21
rect 324 -41 326 -21
rect 499 -36 501 -16
rect 513 -36 515 -16
rect 537 -36 539 -16
rect 561 -36 563 -16
rect 575 -36 577 -16
rect 599 -36 601 -16
rect 623 -36 625 -16
rect 637 -36 639 -16
rect 661 -36 663 -16
rect 1497 -21 1499 -11
rect 1512 -21 1514 -11
rect 1528 -21 1530 -11
rect 1559 -21 1561 -11
rect 1590 -21 1592 -11
rect 11 -98 13 -88
rect 26 -98 28 -88
rect 42 -98 44 -88
rect 73 -98 75 -88
rect 104 -98 106 -88
rect 264 -124 266 -104
rect 1236 -47 1238 -27
rect 1260 -47 1262 -27
rect 1274 -47 1276 -27
rect 1282 -47 1284 -27
rect 1296 -47 1298 -27
rect 499 -133 501 -113
rect 513 -133 515 -113
rect 537 -133 539 -113
rect 561 -133 563 -113
rect 575 -133 577 -113
rect 599 -133 601 -113
rect 729 -120 731 -100
rect 743 -120 745 -100
rect 767 -120 769 -100
rect 791 -120 793 -100
rect 805 -120 807 -100
rect 829 -120 831 -100
rect 853 -120 855 -100
rect 867 -120 869 -100
rect 891 -120 893 -100
rect 1236 -130 1238 -110
rect 1497 -95 1499 -85
rect 1512 -95 1514 -85
rect 1528 -95 1530 -85
rect 1559 -95 1561 -85
rect 1590 -95 1592 -85
rect 11 -172 13 -162
rect 26 -172 28 -162
rect 42 -172 44 -162
rect 73 -172 75 -162
rect 104 -172 106 -162
rect 1497 -169 1499 -159
rect 1512 -169 1514 -159
rect 1528 -169 1530 -159
rect 1559 -169 1561 -159
rect 1590 -169 1592 -159
rect 254 -191 256 -171
rect 268 -191 270 -171
rect 292 -191 294 -171
rect 1236 -197 1238 -177
rect 1260 -197 1262 -177
rect 1274 -197 1276 -177
rect 1282 -197 1284 -177
rect 1296 -197 1298 -177
rect 499 -218 501 -198
rect 513 -218 515 -198
rect 537 -218 539 -198
rect 11 -246 13 -236
rect 26 -246 28 -236
rect 42 -246 44 -236
rect 73 -246 75 -236
rect 104 -246 106 -236
rect 264 -265 266 -245
rect 288 -265 290 -245
rect 302 -265 304 -245
rect 310 -265 312 -245
rect 324 -265 326 -245
rect 11 -320 13 -310
rect 26 -320 28 -310
rect 42 -320 44 -310
rect 73 -320 75 -310
rect 104 -320 106 -310
rect 264 -348 266 -328
rect 1236 -280 1238 -260
rect 1497 -243 1499 -233
rect 1512 -243 1514 -233
rect 1528 -243 1530 -233
rect 1559 -243 1561 -233
rect 1590 -243 1592 -233
rect 499 -330 501 -310
rect 513 -330 515 -310
rect 537 -330 539 -310
rect 561 -330 563 -310
rect 575 -330 577 -310
rect 599 -330 601 -310
rect 623 -330 625 -310
rect 637 -330 639 -310
rect 661 -330 663 -310
rect 685 -330 687 -310
rect 699 -330 701 -310
rect 723 -330 725 -310
rect 1497 -317 1499 -307
rect 1512 -317 1514 -307
rect 1528 -317 1530 -307
rect 1559 -317 1561 -307
rect 1590 -317 1592 -307
rect 1236 -347 1238 -327
rect 1260 -347 1262 -327
rect 1274 -347 1276 -327
rect 1282 -347 1284 -327
rect 1296 -347 1298 -327
rect 11 -394 13 -384
rect 26 -394 28 -384
rect 42 -394 44 -384
rect 73 -394 75 -384
rect 104 -394 106 -384
rect 254 -415 256 -395
rect 268 -415 270 -395
rect 292 -415 294 -395
rect 499 -430 501 -410
rect 513 -430 515 -410
rect 537 -430 539 -410
rect 561 -430 563 -410
rect 575 -430 577 -410
rect 599 -430 601 -410
rect 623 -430 625 -410
rect 637 -430 639 -410
rect 661 -430 663 -410
rect 1236 -430 1238 -410
rect 11 -468 13 -458
rect 26 -468 28 -458
rect 42 -468 44 -458
rect 73 -468 75 -458
rect 104 -468 106 -458
rect 264 -489 266 -469
rect 288 -489 290 -469
rect 302 -489 304 -469
rect 310 -489 312 -469
rect 324 -489 326 -469
rect 264 -572 266 -552
rect 499 -530 501 -510
rect 513 -530 515 -510
rect 537 -530 539 -510
rect 561 -530 563 -510
rect 575 -530 577 -510
rect 599 -530 601 -510
rect 807 -512 809 -492
rect 821 -512 823 -492
rect 845 -512 847 -492
rect 869 -512 871 -492
rect 883 -512 885 -492
rect 907 -512 909 -492
rect 931 -512 933 -492
rect 945 -512 947 -492
rect 969 -512 971 -492
rect 993 -512 995 -492
rect 1007 -512 1009 -492
rect 1031 -512 1033 -492
rect 254 -639 256 -619
rect 268 -639 270 -619
rect 292 -639 294 -619
rect 499 -630 501 -610
rect 513 -630 515 -610
rect 537 -630 539 -610
<< ndiffusion >>
rect 498 195 499 205
rect 501 195 513 205
rect 515 195 516 205
rect 536 195 537 205
rect 539 195 540 205
rect 560 189 561 199
rect 563 189 567 199
rect 571 189 575 199
rect 577 189 578 199
rect 598 189 599 199
rect 601 189 602 199
rect 263 158 264 168
rect 266 158 267 168
rect 498 106 499 116
rect 501 106 513 116
rect 515 106 516 116
rect 536 106 537 116
rect 539 106 540 116
rect 560 106 561 116
rect 563 106 575 116
rect 577 106 578 116
rect 598 106 599 116
rect 601 106 602 116
rect 263 75 264 85
rect 266 75 267 85
rect 287 75 288 85
rect 290 75 291 85
rect 304 75 305 85
rect 307 75 310 85
rect 314 75 318 85
rect 320 75 321 85
rect 334 75 335 85
rect 337 75 338 85
rect 1235 78 1236 88
rect 1238 78 1239 88
rect 641 54 642 64
rect 644 54 648 64
rect 652 54 656 64
rect 658 54 659 64
rect 679 54 680 64
rect 682 54 683 64
rect 703 54 704 64
rect 706 54 710 64
rect 714 54 718 64
rect 720 54 721 64
rect 741 54 742 64
rect 744 54 745 64
rect 10 10 11 20
rect 13 10 14 20
rect 41 10 42 20
rect 44 10 57 20
rect 59 10 60 20
rect 72 10 73 20
rect 75 10 88 20
rect 90 10 91 20
rect 103 10 104 20
rect 106 10 107 20
rect 498 23 499 33
rect 501 23 513 33
rect 515 23 516 33
rect 536 23 537 33
rect 539 23 540 33
rect 253 1 254 11
rect 256 1 268 11
rect 270 1 271 11
rect 291 1 292 11
rect 294 1 295 11
rect 1235 -5 1236 5
rect 1238 -5 1239 5
rect 1259 -5 1260 5
rect 1262 -5 1263 5
rect 1276 -5 1277 5
rect 1279 -5 1282 5
rect 1286 -5 1290 5
rect 1292 -5 1293 5
rect 1306 -5 1307 5
rect 1309 -5 1310 5
rect 10 -64 11 -54
rect 13 -64 14 -54
rect 41 -64 42 -54
rect 44 -64 57 -54
rect 59 -64 60 -54
rect 72 -64 73 -54
rect 75 -64 88 -54
rect 90 -64 91 -54
rect 103 -64 104 -54
rect 106 -64 107 -54
rect 263 -66 264 -56
rect 266 -66 267 -56
rect 10 -138 11 -128
rect 13 -138 14 -128
rect 41 -138 42 -128
rect 44 -138 57 -128
rect 59 -138 60 -128
rect 72 -138 73 -128
rect 75 -138 88 -128
rect 90 -138 91 -128
rect 103 -138 104 -128
rect 106 -138 107 -128
rect 498 -68 499 -58
rect 501 -68 513 -58
rect 515 -68 516 -58
rect 536 -68 537 -58
rect 539 -68 540 -58
rect 560 -68 561 -58
rect 563 -68 575 -58
rect 577 -68 578 -58
rect 598 -68 599 -58
rect 601 -68 602 -58
rect 622 -68 623 -58
rect 625 -68 637 -58
rect 639 -68 640 -58
rect 660 -68 661 -58
rect 663 -68 664 -58
rect 1235 -72 1236 -62
rect 1238 -72 1239 -62
rect 263 -149 264 -139
rect 266 -149 267 -139
rect 287 -149 288 -139
rect 290 -149 291 -139
rect 304 -149 305 -139
rect 307 -149 310 -139
rect 314 -149 318 -139
rect 320 -149 321 -139
rect 334 -149 335 -139
rect 337 -149 338 -139
rect 1496 -61 1497 -51
rect 1499 -61 1500 -51
rect 1527 -61 1528 -51
rect 1530 -61 1543 -51
rect 1545 -61 1546 -51
rect 1558 -61 1559 -51
rect 1561 -61 1574 -51
rect 1576 -61 1577 -51
rect 1589 -61 1590 -51
rect 1592 -61 1593 -51
rect 1496 -135 1497 -125
rect 1499 -135 1500 -125
rect 1527 -135 1528 -125
rect 1530 -135 1543 -125
rect 1545 -135 1546 -125
rect 1558 -135 1559 -125
rect 1561 -135 1574 -125
rect 1576 -135 1577 -125
rect 1589 -135 1590 -125
rect 1592 -135 1593 -125
rect 498 -165 499 -155
rect 501 -165 513 -155
rect 515 -165 516 -155
rect 536 -165 537 -155
rect 539 -165 540 -155
rect 560 -165 561 -155
rect 563 -165 575 -155
rect 577 -165 578 -155
rect 598 -165 599 -155
rect 601 -165 602 -155
rect 728 -158 729 -148
rect 731 -158 735 -148
rect 739 -158 743 -148
rect 745 -158 746 -148
rect 766 -158 767 -148
rect 769 -158 770 -148
rect 790 -158 791 -148
rect 793 -158 797 -148
rect 801 -158 805 -148
rect 807 -158 808 -148
rect 828 -158 829 -148
rect 831 -158 832 -148
rect 852 -158 853 -148
rect 855 -158 859 -148
rect 863 -158 867 -148
rect 869 -158 870 -148
rect 890 -158 891 -148
rect 893 -158 894 -148
rect 1235 -155 1236 -145
rect 1238 -155 1239 -145
rect 1259 -155 1260 -145
rect 1262 -155 1263 -145
rect 1276 -155 1277 -145
rect 1279 -155 1282 -145
rect 1286 -155 1290 -145
rect 1292 -155 1293 -145
rect 1306 -155 1307 -145
rect 1309 -155 1310 -145
rect 10 -212 11 -202
rect 13 -212 14 -202
rect 41 -212 42 -202
rect 44 -212 57 -202
rect 59 -212 60 -202
rect 72 -212 73 -202
rect 75 -212 88 -202
rect 90 -212 91 -202
rect 103 -212 104 -202
rect 106 -212 107 -202
rect 253 -223 254 -213
rect 256 -223 268 -213
rect 270 -223 271 -213
rect 291 -223 292 -213
rect 294 -223 295 -213
rect 1235 -222 1236 -212
rect 1238 -222 1239 -212
rect 498 -250 499 -240
rect 501 -250 513 -240
rect 515 -250 516 -240
rect 536 -250 537 -240
rect 539 -250 540 -240
rect 10 -286 11 -276
rect 13 -286 14 -276
rect 41 -286 42 -276
rect 44 -286 57 -276
rect 59 -286 60 -276
rect 72 -286 73 -276
rect 75 -286 88 -276
rect 90 -286 91 -276
rect 103 -286 104 -276
rect 106 -286 107 -276
rect 263 -290 264 -280
rect 266 -290 267 -280
rect 10 -360 11 -350
rect 13 -360 14 -350
rect 41 -360 42 -350
rect 44 -360 57 -350
rect 59 -360 60 -350
rect 72 -360 73 -350
rect 75 -360 88 -350
rect 90 -360 91 -350
rect 103 -360 104 -350
rect 106 -360 107 -350
rect 1496 -209 1497 -199
rect 1499 -209 1500 -199
rect 1527 -209 1528 -199
rect 1530 -209 1543 -199
rect 1545 -209 1546 -199
rect 1558 -209 1559 -199
rect 1561 -209 1574 -199
rect 1576 -209 1577 -199
rect 1589 -209 1590 -199
rect 1592 -209 1593 -199
rect 1496 -283 1497 -273
rect 1499 -283 1500 -273
rect 1527 -283 1528 -273
rect 1530 -283 1543 -273
rect 1545 -283 1546 -273
rect 1558 -283 1559 -273
rect 1561 -283 1574 -273
rect 1576 -283 1577 -273
rect 1589 -283 1590 -273
rect 1592 -283 1593 -273
rect 1235 -305 1236 -295
rect 1238 -305 1239 -295
rect 1259 -305 1260 -295
rect 1262 -305 1263 -295
rect 1276 -305 1277 -295
rect 1279 -305 1282 -295
rect 1286 -305 1290 -295
rect 1292 -305 1293 -295
rect 1306 -305 1307 -295
rect 1309 -305 1310 -295
rect 498 -362 499 -352
rect 501 -362 513 -352
rect 515 -362 516 -352
rect 536 -362 537 -352
rect 539 -362 540 -352
rect 560 -362 561 -352
rect 563 -362 575 -352
rect 577 -362 578 -352
rect 598 -362 599 -352
rect 601 -362 602 -352
rect 622 -362 623 -352
rect 625 -362 637 -352
rect 639 -362 640 -352
rect 660 -362 661 -352
rect 663 -362 664 -352
rect 684 -362 685 -352
rect 687 -362 699 -352
rect 701 -362 702 -352
rect 722 -362 723 -352
rect 725 -362 726 -352
rect 263 -373 264 -363
rect 266 -373 267 -363
rect 287 -373 288 -363
rect 290 -373 291 -363
rect 304 -373 305 -363
rect 307 -373 310 -363
rect 314 -373 318 -363
rect 320 -373 321 -363
rect 334 -373 335 -363
rect 337 -373 338 -363
rect 1235 -372 1236 -362
rect 1238 -372 1239 -362
rect 10 -434 11 -424
rect 13 -434 14 -424
rect 41 -434 42 -424
rect 44 -434 57 -424
rect 59 -434 60 -424
rect 72 -434 73 -424
rect 75 -434 88 -424
rect 90 -434 91 -424
rect 103 -434 104 -424
rect 106 -434 107 -424
rect 253 -447 254 -437
rect 256 -447 268 -437
rect 270 -447 271 -437
rect 291 -447 292 -437
rect 294 -447 295 -437
rect 1496 -357 1497 -347
rect 1499 -357 1500 -347
rect 1527 -357 1528 -347
rect 1530 -357 1543 -347
rect 1545 -357 1546 -347
rect 1558 -357 1559 -347
rect 1561 -357 1574 -347
rect 1576 -357 1577 -347
rect 1589 -357 1590 -347
rect 1592 -357 1593 -347
rect 498 -462 499 -452
rect 501 -462 513 -452
rect 515 -462 516 -452
rect 536 -462 537 -452
rect 539 -462 540 -452
rect 560 -462 561 -452
rect 563 -462 575 -452
rect 577 -462 578 -452
rect 598 -462 599 -452
rect 601 -462 602 -452
rect 622 -462 623 -452
rect 625 -462 637 -452
rect 639 -462 640 -452
rect 660 -462 661 -452
rect 663 -462 664 -452
rect 1235 -455 1236 -445
rect 1238 -455 1239 -445
rect 1259 -455 1260 -445
rect 1262 -455 1263 -445
rect 1276 -455 1277 -445
rect 1279 -455 1282 -445
rect 1286 -455 1290 -445
rect 1292 -455 1293 -445
rect 1306 -455 1307 -445
rect 1309 -455 1310 -445
rect 10 -508 11 -498
rect 13 -508 14 -498
rect 41 -508 42 -498
rect 44 -508 57 -498
rect 59 -508 60 -498
rect 72 -508 73 -498
rect 75 -508 88 -498
rect 90 -508 91 -498
rect 103 -508 104 -498
rect 106 -508 107 -498
rect 263 -514 264 -504
rect 266 -514 267 -504
rect 806 -550 807 -540
rect 809 -550 813 -540
rect 817 -550 821 -540
rect 823 -550 824 -540
rect 844 -550 845 -540
rect 847 -550 848 -540
rect 868 -550 869 -540
rect 871 -550 875 -540
rect 879 -550 883 -540
rect 885 -550 886 -540
rect 906 -550 907 -540
rect 909 -550 910 -540
rect 930 -550 931 -540
rect 933 -550 937 -540
rect 941 -550 945 -540
rect 947 -550 948 -540
rect 968 -550 969 -540
rect 971 -550 972 -540
rect 992 -550 993 -540
rect 995 -550 999 -540
rect 1003 -550 1007 -540
rect 1009 -550 1010 -540
rect 1030 -550 1031 -540
rect 1033 -550 1034 -540
rect 498 -562 499 -552
rect 501 -562 513 -552
rect 515 -562 516 -552
rect 536 -562 537 -552
rect 539 -562 540 -552
rect 560 -562 561 -552
rect 563 -562 575 -552
rect 577 -562 578 -552
rect 598 -562 599 -552
rect 601 -562 602 -552
rect 263 -597 264 -587
rect 266 -597 267 -587
rect 287 -597 288 -587
rect 290 -597 291 -587
rect 304 -597 305 -587
rect 307 -597 310 -587
rect 314 -597 318 -587
rect 320 -597 321 -587
rect 334 -597 335 -587
rect 337 -597 338 -587
rect 253 -671 254 -661
rect 256 -671 268 -661
rect 270 -671 271 -661
rect 291 -671 292 -661
rect 294 -671 295 -661
rect 498 -662 499 -652
rect 501 -662 513 -652
rect 515 -662 516 -652
rect 536 -662 537 -652
rect 539 -662 540 -652
<< pdiffusion >>
rect 498 227 499 247
rect 501 227 505 247
rect 509 227 513 247
rect 515 227 516 247
rect 536 227 537 247
rect 539 227 540 247
rect 560 227 561 247
rect 563 227 575 247
rect 577 227 578 247
rect 598 227 599 247
rect 601 227 602 247
rect 263 183 264 203
rect 266 183 267 203
rect 287 183 288 203
rect 290 183 302 203
rect 304 183 305 203
rect 309 183 310 203
rect 312 183 324 203
rect 326 183 327 203
rect 263 100 264 120
rect 266 100 267 120
rect 498 138 499 158
rect 501 138 505 158
rect 509 138 513 158
rect 515 138 516 158
rect 536 138 537 158
rect 539 138 540 158
rect 560 138 561 158
rect 563 138 567 158
rect 571 138 575 158
rect 577 138 578 158
rect 598 138 599 158
rect 601 138 602 158
rect 641 92 642 112
rect 644 92 656 112
rect 658 92 659 112
rect 679 92 680 112
rect 682 92 683 112
rect 703 92 704 112
rect 706 92 718 112
rect 720 92 721 112
rect 741 92 742 112
rect 744 92 745 112
rect 1235 103 1236 123
rect 1238 103 1239 123
rect 1259 103 1260 123
rect 1262 103 1274 123
rect 1276 103 1277 123
rect 1281 103 1282 123
rect 1284 103 1296 123
rect 1298 103 1299 123
rect 10 50 11 60
rect 13 50 26 60
rect 28 50 29 60
rect 41 50 42 60
rect 44 50 45 60
rect 72 50 73 60
rect 75 50 76 60
rect 103 50 104 60
rect 106 50 107 60
rect 498 55 499 75
rect 501 55 505 75
rect 509 55 513 75
rect 515 55 516 75
rect 536 55 537 75
rect 539 55 540 75
rect 253 33 254 53
rect 256 33 260 53
rect 264 33 268 53
rect 270 33 271 53
rect 291 33 292 53
rect 294 33 295 53
rect 1235 20 1236 40
rect 1238 20 1239 40
rect 10 -24 11 -14
rect 13 -24 26 -14
rect 28 -24 29 -14
rect 41 -24 42 -14
rect 44 -24 45 -14
rect 72 -24 73 -14
rect 75 -24 76 -14
rect 103 -24 104 -14
rect 106 -24 107 -14
rect 263 -41 264 -21
rect 266 -41 267 -21
rect 287 -41 288 -21
rect 290 -41 302 -21
rect 304 -41 305 -21
rect 309 -41 310 -21
rect 312 -41 324 -21
rect 326 -41 327 -21
rect 498 -36 499 -16
rect 501 -36 505 -16
rect 509 -36 513 -16
rect 515 -36 516 -16
rect 536 -36 537 -16
rect 539 -36 540 -16
rect 560 -36 561 -16
rect 563 -36 567 -16
rect 571 -36 575 -16
rect 577 -36 578 -16
rect 598 -36 599 -16
rect 601 -36 602 -16
rect 622 -36 623 -16
rect 625 -36 629 -16
rect 633 -36 637 -16
rect 639 -36 640 -16
rect 660 -36 661 -16
rect 663 -36 664 -16
rect 1496 -21 1497 -11
rect 1499 -21 1512 -11
rect 1514 -21 1515 -11
rect 1527 -21 1528 -11
rect 1530 -21 1531 -11
rect 1558 -21 1559 -11
rect 1561 -21 1562 -11
rect 1589 -21 1590 -11
rect 1592 -21 1593 -11
rect 10 -98 11 -88
rect 13 -98 26 -88
rect 28 -98 29 -88
rect 41 -98 42 -88
rect 44 -98 45 -88
rect 72 -98 73 -88
rect 75 -98 76 -88
rect 103 -98 104 -88
rect 106 -98 107 -88
rect 263 -124 264 -104
rect 266 -124 267 -104
rect 1235 -47 1236 -27
rect 1238 -47 1239 -27
rect 1259 -47 1260 -27
rect 1262 -47 1274 -27
rect 1276 -47 1277 -27
rect 1281 -47 1282 -27
rect 1284 -47 1296 -27
rect 1298 -47 1299 -27
rect 498 -133 499 -113
rect 501 -133 505 -113
rect 509 -133 513 -113
rect 515 -133 516 -113
rect 536 -133 537 -113
rect 539 -133 540 -113
rect 560 -133 561 -113
rect 563 -133 567 -113
rect 571 -133 575 -113
rect 577 -133 578 -113
rect 598 -133 599 -113
rect 601 -133 602 -113
rect 728 -120 729 -100
rect 731 -120 743 -100
rect 745 -120 746 -100
rect 766 -120 767 -100
rect 769 -120 770 -100
rect 790 -120 791 -100
rect 793 -120 805 -100
rect 807 -120 808 -100
rect 828 -120 829 -100
rect 831 -120 832 -100
rect 852 -120 853 -100
rect 855 -120 867 -100
rect 869 -120 870 -100
rect 890 -120 891 -100
rect 893 -120 894 -100
rect 1235 -130 1236 -110
rect 1238 -130 1239 -110
rect 1496 -95 1497 -85
rect 1499 -95 1512 -85
rect 1514 -95 1515 -85
rect 1527 -95 1528 -85
rect 1530 -95 1531 -85
rect 1558 -95 1559 -85
rect 1561 -95 1562 -85
rect 1589 -95 1590 -85
rect 1592 -95 1593 -85
rect 10 -172 11 -162
rect 13 -172 26 -162
rect 28 -172 29 -162
rect 41 -172 42 -162
rect 44 -172 45 -162
rect 72 -172 73 -162
rect 75 -172 76 -162
rect 103 -172 104 -162
rect 106 -172 107 -162
rect 1496 -169 1497 -159
rect 1499 -169 1512 -159
rect 1514 -169 1515 -159
rect 1527 -169 1528 -159
rect 1530 -169 1531 -159
rect 1558 -169 1559 -159
rect 1561 -169 1562 -159
rect 1589 -169 1590 -159
rect 1592 -169 1593 -159
rect 253 -191 254 -171
rect 256 -191 260 -171
rect 264 -191 268 -171
rect 270 -191 271 -171
rect 291 -191 292 -171
rect 294 -191 295 -171
rect 1235 -197 1236 -177
rect 1238 -197 1239 -177
rect 1259 -197 1260 -177
rect 1262 -197 1274 -177
rect 1276 -197 1277 -177
rect 1281 -197 1282 -177
rect 1284 -197 1296 -177
rect 1298 -197 1299 -177
rect 498 -218 499 -198
rect 501 -218 505 -198
rect 509 -218 513 -198
rect 515 -218 516 -198
rect 536 -218 537 -198
rect 539 -218 540 -198
rect 10 -246 11 -236
rect 13 -246 26 -236
rect 28 -246 29 -236
rect 41 -246 42 -236
rect 44 -246 45 -236
rect 72 -246 73 -236
rect 75 -246 76 -236
rect 103 -246 104 -236
rect 106 -246 107 -236
rect 263 -265 264 -245
rect 266 -265 267 -245
rect 287 -265 288 -245
rect 290 -265 302 -245
rect 304 -265 305 -245
rect 309 -265 310 -245
rect 312 -265 324 -245
rect 326 -265 327 -245
rect 10 -320 11 -310
rect 13 -320 26 -310
rect 28 -320 29 -310
rect 41 -320 42 -310
rect 44 -320 45 -310
rect 72 -320 73 -310
rect 75 -320 76 -310
rect 103 -320 104 -310
rect 106 -320 107 -310
rect 263 -348 264 -328
rect 266 -348 267 -328
rect 1235 -280 1236 -260
rect 1238 -280 1239 -260
rect 1496 -243 1497 -233
rect 1499 -243 1512 -233
rect 1514 -243 1515 -233
rect 1527 -243 1528 -233
rect 1530 -243 1531 -233
rect 1558 -243 1559 -233
rect 1561 -243 1562 -233
rect 1589 -243 1590 -233
rect 1592 -243 1593 -233
rect 498 -330 499 -310
rect 501 -330 505 -310
rect 509 -330 513 -310
rect 515 -330 516 -310
rect 536 -330 537 -310
rect 539 -330 540 -310
rect 560 -330 561 -310
rect 563 -330 567 -310
rect 571 -330 575 -310
rect 577 -330 578 -310
rect 598 -330 599 -310
rect 601 -330 602 -310
rect 622 -330 623 -310
rect 625 -330 629 -310
rect 633 -330 637 -310
rect 639 -330 640 -310
rect 660 -330 661 -310
rect 663 -330 664 -310
rect 684 -330 685 -310
rect 687 -330 691 -310
rect 695 -330 699 -310
rect 701 -330 702 -310
rect 722 -330 723 -310
rect 725 -330 726 -310
rect 1496 -317 1497 -307
rect 1499 -317 1512 -307
rect 1514 -317 1515 -307
rect 1527 -317 1528 -307
rect 1530 -317 1531 -307
rect 1558 -317 1559 -307
rect 1561 -317 1562 -307
rect 1589 -317 1590 -307
rect 1592 -317 1593 -307
rect 1235 -347 1236 -327
rect 1238 -347 1239 -327
rect 1259 -347 1260 -327
rect 1262 -347 1274 -327
rect 1276 -347 1277 -327
rect 1281 -347 1282 -327
rect 1284 -347 1296 -327
rect 1298 -347 1299 -327
rect 10 -394 11 -384
rect 13 -394 26 -384
rect 28 -394 29 -384
rect 41 -394 42 -384
rect 44 -394 45 -384
rect 72 -394 73 -384
rect 75 -394 76 -384
rect 103 -394 104 -384
rect 106 -394 107 -384
rect 253 -415 254 -395
rect 256 -415 260 -395
rect 264 -415 268 -395
rect 270 -415 271 -395
rect 291 -415 292 -395
rect 294 -415 295 -395
rect 498 -430 499 -410
rect 501 -430 505 -410
rect 509 -430 513 -410
rect 515 -430 516 -410
rect 536 -430 537 -410
rect 539 -430 540 -410
rect 560 -430 561 -410
rect 563 -430 567 -410
rect 571 -430 575 -410
rect 577 -430 578 -410
rect 598 -430 599 -410
rect 601 -430 602 -410
rect 622 -430 623 -410
rect 625 -430 629 -410
rect 633 -430 637 -410
rect 639 -430 640 -410
rect 660 -430 661 -410
rect 663 -430 664 -410
rect 1235 -430 1236 -410
rect 1238 -430 1239 -410
rect 10 -468 11 -458
rect 13 -468 26 -458
rect 28 -468 29 -458
rect 41 -468 42 -458
rect 44 -468 45 -458
rect 72 -468 73 -458
rect 75 -468 76 -458
rect 103 -468 104 -458
rect 106 -468 107 -458
rect 263 -489 264 -469
rect 266 -489 267 -469
rect 287 -489 288 -469
rect 290 -489 302 -469
rect 304 -489 305 -469
rect 309 -489 310 -469
rect 312 -489 324 -469
rect 326 -489 327 -469
rect 263 -572 264 -552
rect 266 -572 267 -552
rect 498 -530 499 -510
rect 501 -530 505 -510
rect 509 -530 513 -510
rect 515 -530 516 -510
rect 536 -530 537 -510
rect 539 -530 540 -510
rect 560 -530 561 -510
rect 563 -530 567 -510
rect 571 -530 575 -510
rect 577 -530 578 -510
rect 598 -530 599 -510
rect 601 -530 602 -510
rect 806 -512 807 -492
rect 809 -512 821 -492
rect 823 -512 824 -492
rect 844 -512 845 -492
rect 847 -512 848 -492
rect 868 -512 869 -492
rect 871 -512 883 -492
rect 885 -512 886 -492
rect 906 -512 907 -492
rect 909 -512 910 -492
rect 930 -512 931 -492
rect 933 -512 945 -492
rect 947 -512 948 -492
rect 968 -512 969 -492
rect 971 -512 972 -492
rect 992 -512 993 -492
rect 995 -512 1007 -492
rect 1009 -512 1010 -492
rect 1030 -512 1031 -492
rect 1033 -512 1034 -492
rect 253 -639 254 -619
rect 256 -639 260 -619
rect 264 -639 268 -619
rect 270 -639 271 -619
rect 291 -639 292 -619
rect 294 -639 295 -619
rect 498 -630 499 -610
rect 501 -630 505 -610
rect 509 -630 513 -610
rect 515 -630 516 -610
rect 536 -630 537 -610
rect 539 -630 540 -610
<< ndcontact >>
rect 494 195 498 205
rect 516 195 520 205
rect 532 195 536 205
rect 540 195 544 205
rect 556 189 560 199
rect 567 189 571 199
rect 578 189 582 199
rect 594 189 598 199
rect 602 189 606 199
rect 259 158 263 168
rect 267 158 271 168
rect 494 106 498 116
rect 516 106 520 116
rect 532 106 536 116
rect 540 106 544 116
rect 556 106 560 116
rect 578 106 582 116
rect 594 106 598 116
rect 602 106 606 116
rect 259 75 263 85
rect 267 75 271 85
rect 283 75 287 85
rect 291 75 295 85
rect 310 75 314 85
rect 321 75 325 85
rect 338 75 342 85
rect 1231 78 1235 88
rect 1239 78 1243 88
rect 637 54 641 64
rect 648 54 652 64
rect 659 54 663 64
rect 675 54 679 64
rect 683 54 687 64
rect 699 54 703 64
rect 710 54 714 64
rect 721 54 725 64
rect 737 54 741 64
rect 745 54 749 64
rect 6 10 10 20
rect 14 10 18 20
rect 37 10 41 20
rect 60 10 64 20
rect 68 10 72 20
rect 91 10 95 20
rect 99 10 103 20
rect 107 10 111 20
rect 494 23 498 33
rect 516 23 520 33
rect 532 23 536 33
rect 540 23 544 33
rect 249 1 253 11
rect 271 1 275 11
rect 287 1 291 11
rect 295 1 299 11
rect 1231 -5 1235 5
rect 1239 -5 1243 5
rect 1255 -5 1259 5
rect 1263 -5 1267 5
rect 1282 -5 1286 5
rect 1293 -5 1297 5
rect 1310 -5 1314 5
rect 6 -64 10 -54
rect 14 -64 18 -54
rect 37 -64 41 -54
rect 60 -64 64 -54
rect 68 -64 72 -54
rect 91 -64 95 -54
rect 99 -64 103 -54
rect 107 -64 111 -54
rect 259 -66 263 -56
rect 267 -66 271 -56
rect 6 -138 10 -128
rect 14 -138 18 -128
rect 37 -138 41 -128
rect 60 -138 64 -128
rect 68 -138 72 -128
rect 91 -138 95 -128
rect 99 -138 103 -128
rect 107 -138 111 -128
rect 494 -68 498 -58
rect 516 -68 520 -58
rect 532 -68 536 -58
rect 540 -68 544 -58
rect 556 -68 560 -58
rect 578 -68 582 -58
rect 594 -68 598 -58
rect 602 -68 606 -58
rect 618 -68 622 -58
rect 640 -68 644 -58
rect 656 -68 660 -58
rect 664 -68 668 -58
rect 1231 -72 1235 -62
rect 1239 -72 1243 -62
rect 259 -149 263 -139
rect 267 -149 271 -139
rect 283 -149 287 -139
rect 291 -149 295 -139
rect 310 -149 314 -139
rect 321 -149 325 -139
rect 338 -149 342 -139
rect 1492 -61 1496 -51
rect 1500 -61 1504 -51
rect 1523 -61 1527 -51
rect 1546 -61 1550 -51
rect 1554 -61 1558 -51
rect 1577 -61 1581 -51
rect 1585 -61 1589 -51
rect 1593 -61 1597 -51
rect 1492 -135 1496 -125
rect 1500 -135 1504 -125
rect 1523 -135 1527 -125
rect 1546 -135 1550 -125
rect 1554 -135 1558 -125
rect 1577 -135 1581 -125
rect 1585 -135 1589 -125
rect 1593 -135 1597 -125
rect 494 -165 498 -155
rect 516 -165 520 -155
rect 532 -165 536 -155
rect 540 -165 544 -155
rect 556 -165 560 -155
rect 578 -165 582 -155
rect 594 -165 598 -155
rect 602 -165 606 -155
rect 724 -158 728 -148
rect 735 -158 739 -148
rect 746 -158 750 -148
rect 762 -158 766 -148
rect 770 -158 774 -148
rect 786 -158 790 -148
rect 797 -158 801 -148
rect 808 -158 812 -148
rect 824 -158 828 -148
rect 832 -158 836 -148
rect 848 -158 852 -148
rect 859 -158 863 -148
rect 870 -158 874 -148
rect 886 -158 890 -148
rect 894 -158 898 -148
rect 1231 -155 1235 -145
rect 1239 -155 1243 -145
rect 1255 -155 1259 -145
rect 1263 -155 1267 -145
rect 1282 -155 1286 -145
rect 1293 -155 1297 -145
rect 1310 -155 1314 -145
rect 6 -212 10 -202
rect 14 -212 18 -202
rect 37 -212 41 -202
rect 60 -212 64 -202
rect 68 -212 72 -202
rect 91 -212 95 -202
rect 99 -212 103 -202
rect 107 -212 111 -202
rect 249 -223 253 -213
rect 271 -223 275 -213
rect 287 -223 291 -213
rect 295 -223 299 -213
rect 1231 -222 1235 -212
rect 1239 -222 1243 -212
rect 494 -250 498 -240
rect 516 -250 520 -240
rect 532 -250 536 -240
rect 540 -250 544 -240
rect 6 -286 10 -276
rect 14 -286 18 -276
rect 37 -286 41 -276
rect 60 -286 64 -276
rect 68 -286 72 -276
rect 91 -286 95 -276
rect 99 -286 103 -276
rect 107 -286 111 -276
rect 259 -290 263 -280
rect 267 -290 271 -280
rect 6 -360 10 -350
rect 14 -360 18 -350
rect 37 -360 41 -350
rect 60 -360 64 -350
rect 68 -360 72 -350
rect 91 -360 95 -350
rect 99 -360 103 -350
rect 107 -360 111 -350
rect 1492 -209 1496 -199
rect 1500 -209 1504 -199
rect 1523 -209 1527 -199
rect 1546 -209 1550 -199
rect 1554 -209 1558 -199
rect 1577 -209 1581 -199
rect 1585 -209 1589 -199
rect 1593 -209 1597 -199
rect 1492 -283 1496 -273
rect 1500 -283 1504 -273
rect 1523 -283 1527 -273
rect 1546 -283 1550 -273
rect 1554 -283 1558 -273
rect 1577 -283 1581 -273
rect 1585 -283 1589 -273
rect 1593 -283 1597 -273
rect 1231 -305 1235 -295
rect 1239 -305 1243 -295
rect 1255 -305 1259 -295
rect 1263 -305 1267 -295
rect 1282 -305 1286 -295
rect 1293 -305 1297 -295
rect 1310 -305 1314 -295
rect 494 -362 498 -352
rect 516 -362 520 -352
rect 532 -362 536 -352
rect 540 -362 544 -352
rect 556 -362 560 -352
rect 578 -362 582 -352
rect 594 -362 598 -352
rect 602 -362 606 -352
rect 618 -362 622 -352
rect 640 -362 644 -352
rect 656 -362 660 -352
rect 664 -362 668 -352
rect 680 -362 684 -352
rect 702 -362 706 -352
rect 718 -362 722 -352
rect 726 -362 730 -352
rect 259 -373 263 -363
rect 267 -373 271 -363
rect 283 -373 287 -363
rect 291 -373 295 -363
rect 310 -373 314 -363
rect 321 -373 325 -363
rect 338 -373 342 -363
rect 1231 -372 1235 -362
rect 1239 -372 1243 -362
rect 6 -434 10 -424
rect 14 -434 18 -424
rect 37 -434 41 -424
rect 60 -434 64 -424
rect 68 -434 72 -424
rect 91 -434 95 -424
rect 99 -434 103 -424
rect 107 -434 111 -424
rect 249 -447 253 -437
rect 271 -447 275 -437
rect 287 -447 291 -437
rect 295 -447 299 -437
rect 1492 -357 1496 -347
rect 1500 -357 1504 -347
rect 1523 -357 1527 -347
rect 1546 -357 1550 -347
rect 1554 -357 1558 -347
rect 1577 -357 1581 -347
rect 1585 -357 1589 -347
rect 1593 -357 1597 -347
rect 494 -462 498 -452
rect 516 -462 520 -452
rect 532 -462 536 -452
rect 540 -462 544 -452
rect 556 -462 560 -452
rect 578 -462 582 -452
rect 594 -462 598 -452
rect 602 -462 606 -452
rect 618 -462 622 -452
rect 640 -462 644 -452
rect 656 -462 660 -452
rect 664 -462 668 -452
rect 1231 -455 1235 -445
rect 1239 -455 1243 -445
rect 1255 -455 1259 -445
rect 1263 -455 1267 -445
rect 1282 -455 1286 -445
rect 1293 -455 1297 -445
rect 1310 -455 1314 -445
rect 6 -508 10 -498
rect 14 -508 18 -498
rect 37 -508 41 -498
rect 60 -508 64 -498
rect 68 -508 72 -498
rect 91 -508 95 -498
rect 99 -508 103 -498
rect 107 -508 111 -498
rect 259 -514 263 -504
rect 267 -514 271 -504
rect 802 -550 806 -540
rect 813 -550 817 -540
rect 824 -550 828 -540
rect 840 -550 844 -540
rect 848 -550 852 -540
rect 864 -550 868 -540
rect 875 -550 879 -540
rect 886 -550 890 -540
rect 902 -550 906 -540
rect 910 -550 914 -540
rect 926 -550 930 -540
rect 937 -550 941 -540
rect 948 -550 952 -540
rect 964 -550 968 -540
rect 972 -550 976 -540
rect 988 -550 992 -540
rect 999 -550 1003 -540
rect 1010 -550 1014 -540
rect 1026 -550 1030 -540
rect 1034 -550 1038 -540
rect 494 -562 498 -552
rect 516 -562 520 -552
rect 532 -562 536 -552
rect 540 -562 544 -552
rect 556 -562 560 -552
rect 578 -562 582 -552
rect 594 -562 598 -552
rect 602 -562 606 -552
rect 259 -597 263 -587
rect 267 -597 271 -587
rect 283 -597 287 -587
rect 291 -597 295 -587
rect 310 -597 314 -587
rect 321 -597 325 -587
rect 338 -597 342 -587
rect 249 -671 253 -661
rect 271 -671 275 -661
rect 287 -671 291 -661
rect 295 -671 299 -661
rect 494 -662 498 -652
rect 516 -662 520 -652
rect 532 -662 536 -652
rect 540 -662 544 -652
<< pdcontact >>
rect 494 227 498 247
rect 505 227 509 247
rect 516 227 520 247
rect 532 227 536 247
rect 540 227 544 247
rect 556 227 560 247
rect 578 227 582 247
rect 594 227 598 247
rect 602 227 606 247
rect 259 183 263 203
rect 267 183 271 203
rect 283 183 287 203
rect 305 183 309 203
rect 327 183 331 203
rect 259 100 263 120
rect 267 100 271 120
rect 494 138 498 158
rect 505 138 509 158
rect 516 138 520 158
rect 532 138 536 158
rect 540 138 544 158
rect 556 138 560 158
rect 567 138 571 158
rect 578 138 582 158
rect 594 138 598 158
rect 602 138 606 158
rect 637 92 641 112
rect 659 92 663 112
rect 675 92 679 112
rect 683 92 687 112
rect 699 92 703 112
rect 721 92 725 112
rect 737 92 741 112
rect 745 92 749 112
rect 1231 103 1235 123
rect 1239 103 1243 123
rect 1255 103 1259 123
rect 1277 103 1281 123
rect 1299 103 1303 123
rect 6 50 10 60
rect 29 50 33 60
rect 37 50 41 60
rect 45 50 49 60
rect 68 50 72 60
rect 76 50 80 60
rect 99 50 103 60
rect 107 50 111 60
rect 494 55 498 75
rect 505 55 509 75
rect 516 55 520 75
rect 532 55 536 75
rect 540 55 544 75
rect 249 33 253 53
rect 260 33 264 53
rect 271 33 275 53
rect 287 33 291 53
rect 295 33 299 53
rect 1231 20 1235 40
rect 1239 20 1243 40
rect 6 -24 10 -14
rect 29 -24 33 -14
rect 37 -24 41 -14
rect 45 -24 49 -14
rect 68 -24 72 -14
rect 76 -24 80 -14
rect 99 -24 103 -14
rect 107 -24 111 -14
rect 259 -41 263 -21
rect 267 -41 271 -21
rect 283 -41 287 -21
rect 305 -41 309 -21
rect 327 -41 331 -21
rect 494 -36 498 -16
rect 505 -36 509 -16
rect 516 -36 520 -16
rect 532 -36 536 -16
rect 540 -36 544 -16
rect 556 -36 560 -16
rect 567 -36 571 -16
rect 578 -36 582 -16
rect 594 -36 598 -16
rect 602 -36 606 -16
rect 618 -36 622 -16
rect 629 -36 633 -16
rect 640 -36 644 -16
rect 656 -36 660 -16
rect 664 -36 668 -16
rect 1492 -21 1496 -11
rect 1515 -21 1519 -11
rect 1523 -21 1527 -11
rect 1531 -21 1535 -11
rect 1554 -21 1558 -11
rect 1562 -21 1566 -11
rect 1585 -21 1589 -11
rect 1593 -21 1597 -11
rect 6 -98 10 -88
rect 29 -98 33 -88
rect 37 -98 41 -88
rect 45 -98 49 -88
rect 68 -98 72 -88
rect 76 -98 80 -88
rect 99 -98 103 -88
rect 107 -98 111 -88
rect 259 -124 263 -104
rect 267 -124 271 -104
rect 1231 -47 1235 -27
rect 1239 -47 1243 -27
rect 1255 -47 1259 -27
rect 1277 -47 1281 -27
rect 1299 -47 1303 -27
rect 494 -133 498 -113
rect 505 -133 509 -113
rect 516 -133 520 -113
rect 532 -133 536 -113
rect 540 -133 544 -113
rect 556 -133 560 -113
rect 567 -133 571 -113
rect 578 -133 582 -113
rect 594 -133 598 -113
rect 602 -133 606 -113
rect 724 -120 728 -100
rect 746 -120 750 -100
rect 762 -120 766 -100
rect 770 -120 774 -100
rect 786 -120 790 -100
rect 808 -120 812 -100
rect 824 -120 828 -100
rect 832 -120 836 -100
rect 848 -120 852 -100
rect 870 -120 874 -100
rect 886 -120 890 -100
rect 894 -120 898 -100
rect 1231 -130 1235 -110
rect 1239 -130 1243 -110
rect 1492 -95 1496 -85
rect 1515 -95 1519 -85
rect 1523 -95 1527 -85
rect 1531 -95 1535 -85
rect 1554 -95 1558 -85
rect 1562 -95 1566 -85
rect 1585 -95 1589 -85
rect 1593 -95 1597 -85
rect 6 -172 10 -162
rect 29 -172 33 -162
rect 37 -172 41 -162
rect 45 -172 49 -162
rect 68 -172 72 -162
rect 76 -172 80 -162
rect 99 -172 103 -162
rect 107 -172 111 -162
rect 1492 -169 1496 -159
rect 1515 -169 1519 -159
rect 1523 -169 1527 -159
rect 1531 -169 1535 -159
rect 1554 -169 1558 -159
rect 1562 -169 1566 -159
rect 1585 -169 1589 -159
rect 1593 -169 1597 -159
rect 249 -191 253 -171
rect 260 -191 264 -171
rect 271 -191 275 -171
rect 287 -191 291 -171
rect 295 -191 299 -171
rect 1231 -197 1235 -177
rect 1239 -197 1243 -177
rect 1255 -197 1259 -177
rect 1277 -197 1281 -177
rect 1299 -197 1303 -177
rect 494 -218 498 -198
rect 505 -218 509 -198
rect 516 -218 520 -198
rect 532 -218 536 -198
rect 540 -218 544 -198
rect 6 -246 10 -236
rect 29 -246 33 -236
rect 37 -246 41 -236
rect 45 -246 49 -236
rect 68 -246 72 -236
rect 76 -246 80 -236
rect 99 -246 103 -236
rect 107 -246 111 -236
rect 259 -265 263 -245
rect 267 -265 271 -245
rect 283 -265 287 -245
rect 305 -265 309 -245
rect 327 -265 331 -245
rect 6 -320 10 -310
rect 29 -320 33 -310
rect 37 -320 41 -310
rect 45 -320 49 -310
rect 68 -320 72 -310
rect 76 -320 80 -310
rect 99 -320 103 -310
rect 107 -320 111 -310
rect 259 -348 263 -328
rect 267 -348 271 -328
rect 1231 -280 1235 -260
rect 1239 -280 1243 -260
rect 1492 -243 1496 -233
rect 1515 -243 1519 -233
rect 1523 -243 1527 -233
rect 1531 -243 1535 -233
rect 1554 -243 1558 -233
rect 1562 -243 1566 -233
rect 1585 -243 1589 -233
rect 1593 -243 1597 -233
rect 494 -330 498 -310
rect 505 -330 509 -310
rect 516 -330 520 -310
rect 532 -330 536 -310
rect 540 -330 544 -310
rect 556 -330 560 -310
rect 567 -330 571 -310
rect 578 -330 582 -310
rect 594 -330 598 -310
rect 602 -330 606 -310
rect 618 -330 622 -310
rect 629 -330 633 -310
rect 640 -330 644 -310
rect 656 -330 660 -310
rect 664 -330 668 -310
rect 680 -330 684 -310
rect 691 -330 695 -310
rect 702 -330 706 -310
rect 718 -330 722 -310
rect 726 -330 730 -310
rect 1492 -317 1496 -307
rect 1515 -317 1519 -307
rect 1523 -317 1527 -307
rect 1531 -317 1535 -307
rect 1554 -317 1558 -307
rect 1562 -317 1566 -307
rect 1585 -317 1589 -307
rect 1593 -317 1597 -307
rect 1231 -347 1235 -327
rect 1239 -347 1243 -327
rect 1255 -347 1259 -327
rect 1277 -347 1281 -327
rect 1299 -347 1303 -327
rect 6 -394 10 -384
rect 29 -394 33 -384
rect 37 -394 41 -384
rect 45 -394 49 -384
rect 68 -394 72 -384
rect 76 -394 80 -384
rect 99 -394 103 -384
rect 107 -394 111 -384
rect 249 -415 253 -395
rect 260 -415 264 -395
rect 271 -415 275 -395
rect 287 -415 291 -395
rect 295 -415 299 -395
rect 494 -430 498 -410
rect 505 -430 509 -410
rect 516 -430 520 -410
rect 532 -430 536 -410
rect 540 -430 544 -410
rect 556 -430 560 -410
rect 567 -430 571 -410
rect 578 -430 582 -410
rect 594 -430 598 -410
rect 602 -430 606 -410
rect 618 -430 622 -410
rect 629 -430 633 -410
rect 640 -430 644 -410
rect 656 -430 660 -410
rect 664 -430 668 -410
rect 1231 -430 1235 -410
rect 1239 -430 1243 -410
rect 6 -468 10 -458
rect 29 -468 33 -458
rect 37 -468 41 -458
rect 45 -468 49 -458
rect 68 -468 72 -458
rect 76 -468 80 -458
rect 99 -468 103 -458
rect 107 -468 111 -458
rect 259 -489 263 -469
rect 267 -489 271 -469
rect 283 -489 287 -469
rect 305 -489 309 -469
rect 327 -489 331 -469
rect 259 -572 263 -552
rect 267 -572 271 -552
rect 494 -530 498 -510
rect 505 -530 509 -510
rect 516 -530 520 -510
rect 532 -530 536 -510
rect 540 -530 544 -510
rect 556 -530 560 -510
rect 567 -530 571 -510
rect 578 -530 582 -510
rect 594 -530 598 -510
rect 602 -530 606 -510
rect 802 -512 806 -492
rect 824 -512 828 -492
rect 840 -512 844 -492
rect 848 -512 852 -492
rect 864 -512 868 -492
rect 886 -512 890 -492
rect 902 -512 906 -492
rect 910 -512 914 -492
rect 926 -512 930 -492
rect 948 -512 952 -492
rect 964 -512 968 -492
rect 972 -512 976 -492
rect 988 -512 992 -492
rect 1010 -512 1014 -492
rect 1026 -512 1030 -492
rect 1034 -512 1038 -492
rect 249 -639 253 -619
rect 260 -639 264 -619
rect 271 -639 275 -619
rect 287 -639 291 -619
rect 295 -639 299 -619
rect 494 -630 498 -610
rect 505 -630 509 -610
rect 516 -630 520 -610
rect 532 -630 536 -610
rect 540 -630 544 -610
<< psubstratepcontact >>
rect 536 187 540 191
rect 598 181 602 185
rect 536 98 540 102
rect 598 98 602 102
rect 263 67 267 71
rect 679 46 683 50
rect 741 46 745 50
rect 536 15 540 19
rect 52 0 56 4
rect 291 -7 295 -3
rect 1235 -13 1239 -9
rect 52 -74 56 -70
rect 536 -76 540 -72
rect 598 -76 602 -72
rect 660 -76 664 -72
rect 52 -148 56 -144
rect 263 -157 267 -153
rect 1538 -71 1542 -67
rect 1538 -145 1542 -141
rect 766 -166 770 -162
rect 828 -166 832 -162
rect 890 -166 894 -162
rect 1235 -163 1239 -159
rect 536 -173 540 -169
rect 598 -173 602 -169
rect 52 -222 56 -218
rect 291 -231 295 -227
rect 536 -258 540 -254
rect 52 -296 56 -292
rect 1538 -219 1542 -215
rect 1538 -293 1542 -289
rect 1235 -313 1239 -309
rect 52 -370 56 -366
rect 536 -370 540 -366
rect 598 -370 602 -366
rect 660 -370 664 -366
rect 722 -370 726 -366
rect 263 -381 267 -377
rect 52 -444 56 -440
rect 291 -455 295 -451
rect 1538 -367 1542 -363
rect 1235 -463 1239 -459
rect 536 -470 540 -466
rect 598 -470 602 -466
rect 660 -470 664 -466
rect 52 -518 56 -514
rect 844 -558 848 -554
rect 906 -558 910 -554
rect 968 -558 972 -554
rect 1030 -558 1034 -554
rect 536 -570 540 -566
rect 598 -570 602 -566
rect 263 -605 267 -601
rect 536 -670 540 -666
rect 291 -679 295 -675
<< nsubstratencontact >>
rect 536 251 540 255
rect 598 251 602 255
rect 263 207 267 211
rect 263 124 267 128
rect 536 162 540 166
rect 598 162 602 166
rect 1235 127 1239 131
rect 679 116 683 120
rect 741 116 745 120
rect 536 79 540 83
rect 54 64 58 68
rect 291 57 295 61
rect 1235 44 1239 48
rect 54 -10 58 -6
rect 1540 -7 1544 -3
rect 536 -12 540 -8
rect 598 -12 602 -8
rect 660 -12 664 -8
rect 263 -17 267 -13
rect 1235 -23 1239 -19
rect 54 -84 58 -80
rect 263 -100 267 -96
rect 766 -96 770 -92
rect 828 -96 832 -92
rect 890 -96 894 -92
rect 536 -109 540 -105
rect 598 -109 602 -105
rect 1235 -106 1239 -102
rect 54 -158 58 -154
rect 1540 -81 1544 -77
rect 291 -167 295 -163
rect 1540 -155 1544 -151
rect 1235 -173 1239 -169
rect 536 -194 540 -190
rect 54 -232 58 -228
rect 263 -241 267 -237
rect 1235 -256 1239 -252
rect 54 -306 58 -302
rect 263 -324 267 -320
rect 1540 -229 1544 -225
rect 536 -306 540 -302
rect 598 -306 602 -302
rect 660 -306 664 -302
rect 722 -306 726 -302
rect 1540 -303 1544 -299
rect 1235 -323 1239 -319
rect 54 -380 58 -376
rect 291 -391 295 -387
rect 536 -406 540 -402
rect 598 -406 602 -402
rect 660 -406 664 -402
rect 1235 -406 1239 -402
rect 54 -454 58 -450
rect 263 -465 267 -461
rect 844 -488 848 -484
rect 906 -488 910 -484
rect 968 -488 972 -484
rect 1030 -488 1034 -484
rect 263 -548 267 -544
rect 536 -506 540 -502
rect 598 -506 602 -502
rect 536 -606 540 -602
rect 291 -615 295 -611
<< polysilicon >>
rect 499 247 501 250
rect 513 247 515 250
rect 537 247 539 250
rect 561 247 563 250
rect 575 247 577 250
rect 599 247 601 250
rect 264 203 266 206
rect 288 203 290 206
rect 302 203 304 206
rect 310 203 312 206
rect 324 203 326 206
rect 499 205 501 227
rect 513 205 515 227
rect 537 205 539 227
rect 561 199 563 227
rect 575 199 577 227
rect 599 199 601 227
rect 499 192 501 195
rect 513 192 515 195
rect 537 192 539 195
rect 561 186 563 189
rect 575 186 577 189
rect 599 186 601 189
rect 264 168 266 183
rect 264 155 266 158
rect 264 120 266 123
rect 264 85 266 100
rect 288 85 290 183
rect 302 112 304 183
rect 297 110 304 112
rect 297 97 299 110
rect 297 95 304 97
rect 302 88 304 95
rect 310 88 312 183
rect 324 88 326 183
rect 499 158 501 161
rect 513 158 515 161
rect 537 158 539 161
rect 561 158 563 161
rect 575 158 577 161
rect 599 158 601 161
rect 499 116 501 138
rect 513 116 515 138
rect 537 116 539 138
rect 561 116 563 138
rect 575 116 577 138
rect 599 116 601 138
rect 1236 123 1238 126
rect 1260 123 1262 126
rect 1274 123 1276 126
rect 1282 123 1284 126
rect 1296 123 1298 126
rect 642 112 644 115
rect 656 112 658 115
rect 680 112 682 115
rect 704 112 706 115
rect 718 112 720 115
rect 742 112 744 115
rect 499 103 501 106
rect 513 103 515 106
rect 537 103 539 106
rect 561 103 563 106
rect 575 103 577 106
rect 599 103 601 106
rect 302 86 307 88
rect 310 86 320 88
rect 324 86 337 88
rect 305 85 307 86
rect 318 85 320 86
rect 335 85 337 86
rect 499 75 501 78
rect 513 75 515 78
rect 537 75 539 78
rect 264 72 266 75
rect 288 72 290 75
rect 305 72 307 75
rect 318 72 320 75
rect 335 72 337 75
rect 11 60 13 63
rect 26 60 28 63
rect 42 60 44 63
rect 73 60 75 63
rect 104 60 106 63
rect 254 53 256 56
rect 268 53 270 56
rect 292 53 294 56
rect 642 64 644 92
rect 656 64 658 92
rect 680 64 682 92
rect 704 64 706 92
rect 718 64 720 92
rect 742 64 744 92
rect 1236 88 1238 103
rect 1236 75 1238 78
rect 11 20 13 50
rect 26 36 28 50
rect 42 20 44 50
rect 57 20 59 32
rect 73 20 75 50
rect 88 20 90 41
rect 104 20 106 50
rect 499 33 501 55
rect 513 33 515 55
rect 537 33 539 55
rect 642 51 644 54
rect 656 51 658 54
rect 680 51 682 54
rect 704 51 706 54
rect 718 51 720 54
rect 742 51 744 54
rect 1236 40 1238 43
rect 254 11 256 33
rect 268 11 270 33
rect 292 11 294 33
rect 499 20 501 23
rect 513 20 515 23
rect 537 20 539 23
rect 11 7 13 10
rect 42 7 44 10
rect 57 7 59 10
rect 73 7 75 10
rect 88 7 90 10
rect 104 7 106 10
rect 1236 5 1238 20
rect 1260 5 1262 103
rect 1274 32 1276 103
rect 1269 30 1276 32
rect 1269 17 1271 30
rect 1269 15 1276 17
rect 1274 8 1276 15
rect 1282 8 1284 103
rect 1296 8 1298 103
rect 1274 6 1279 8
rect 1282 6 1292 8
rect 1296 6 1309 8
rect 1277 5 1279 6
rect 1290 5 1292 6
rect 1307 5 1309 6
rect 254 -2 256 1
rect 268 -2 270 1
rect 292 -2 294 1
rect 1236 -8 1238 -5
rect 1260 -8 1262 -5
rect 1277 -8 1279 -5
rect 1290 -8 1292 -5
rect 1307 -8 1309 -5
rect 11 -14 13 -11
rect 26 -14 28 -11
rect 42 -14 44 -11
rect 73 -14 75 -11
rect 104 -14 106 -11
rect 1497 -11 1499 -8
rect 1512 -11 1514 -8
rect 1528 -11 1530 -8
rect 1559 -11 1561 -8
rect 1590 -11 1592 -8
rect 499 -16 501 -13
rect 513 -16 515 -13
rect 537 -16 539 -13
rect 561 -16 563 -13
rect 575 -16 577 -13
rect 599 -16 601 -13
rect 623 -16 625 -13
rect 637 -16 639 -13
rect 661 -16 663 -13
rect 264 -21 266 -18
rect 288 -21 290 -18
rect 302 -21 304 -18
rect 310 -21 312 -18
rect 324 -21 326 -18
rect 11 -54 13 -24
rect 26 -38 28 -24
rect 42 -54 44 -24
rect 57 -54 59 -42
rect 73 -54 75 -24
rect 88 -54 90 -33
rect 104 -54 106 -24
rect 1236 -27 1238 -24
rect 1260 -27 1262 -24
rect 1274 -27 1276 -24
rect 1282 -27 1284 -24
rect 1296 -27 1298 -24
rect 264 -56 266 -41
rect 11 -67 13 -64
rect 42 -67 44 -64
rect 57 -67 59 -64
rect 73 -67 75 -64
rect 88 -67 90 -64
rect 104 -67 106 -64
rect 264 -69 266 -66
rect 11 -88 13 -85
rect 26 -88 28 -85
rect 42 -88 44 -85
rect 73 -88 75 -85
rect 104 -88 106 -85
rect 11 -128 13 -98
rect 26 -112 28 -98
rect 42 -128 44 -98
rect 57 -128 59 -116
rect 73 -128 75 -98
rect 88 -128 90 -107
rect 104 -128 106 -98
rect 264 -104 266 -101
rect 11 -141 13 -138
rect 42 -141 44 -138
rect 57 -141 59 -138
rect 73 -141 75 -138
rect 88 -141 90 -138
rect 104 -141 106 -138
rect 264 -139 266 -124
rect 288 -139 290 -41
rect 302 -112 304 -41
rect 297 -114 304 -112
rect 297 -127 299 -114
rect 297 -129 304 -127
rect 302 -136 304 -129
rect 310 -136 312 -41
rect 324 -136 326 -41
rect 499 -58 501 -36
rect 513 -58 515 -36
rect 537 -58 539 -36
rect 561 -58 563 -36
rect 575 -58 577 -36
rect 599 -58 601 -36
rect 623 -58 625 -36
rect 637 -58 639 -36
rect 661 -58 663 -36
rect 1236 -62 1238 -47
rect 499 -71 501 -68
rect 513 -71 515 -68
rect 537 -71 539 -68
rect 561 -71 563 -68
rect 575 -71 577 -68
rect 599 -71 601 -68
rect 623 -71 625 -68
rect 637 -71 639 -68
rect 661 -71 663 -68
rect 1236 -75 1238 -72
rect 729 -100 731 -97
rect 743 -100 745 -97
rect 767 -100 769 -97
rect 791 -100 793 -97
rect 805 -100 807 -97
rect 829 -100 831 -97
rect 853 -100 855 -97
rect 867 -100 869 -97
rect 891 -100 893 -97
rect 499 -113 501 -110
rect 513 -113 515 -110
rect 537 -113 539 -110
rect 561 -113 563 -110
rect 575 -113 577 -110
rect 599 -113 601 -110
rect 1236 -110 1238 -107
rect 302 -138 307 -136
rect 310 -138 320 -136
rect 324 -138 337 -136
rect 305 -139 307 -138
rect 318 -139 320 -138
rect 335 -139 337 -138
rect 264 -152 266 -149
rect 288 -152 290 -149
rect 305 -152 307 -149
rect 318 -152 320 -149
rect 335 -152 337 -149
rect 499 -155 501 -133
rect 513 -155 515 -133
rect 537 -155 539 -133
rect 561 -155 563 -133
rect 575 -155 577 -133
rect 599 -155 601 -133
rect 729 -148 731 -120
rect 743 -148 745 -120
rect 767 -148 769 -120
rect 791 -148 793 -120
rect 805 -148 807 -120
rect 829 -148 831 -120
rect 853 -148 855 -120
rect 867 -148 869 -120
rect 891 -148 893 -120
rect 1236 -145 1238 -130
rect 1260 -145 1262 -47
rect 1274 -118 1276 -47
rect 1269 -120 1276 -118
rect 1269 -133 1271 -120
rect 1269 -135 1276 -133
rect 1274 -142 1276 -135
rect 1282 -142 1284 -47
rect 1296 -142 1298 -47
rect 1497 -51 1499 -21
rect 1512 -35 1514 -21
rect 1528 -51 1530 -21
rect 1543 -51 1545 -39
rect 1559 -51 1561 -21
rect 1574 -51 1576 -30
rect 1590 -51 1592 -21
rect 1497 -64 1499 -61
rect 1528 -64 1530 -61
rect 1543 -64 1545 -61
rect 1559 -64 1561 -61
rect 1574 -64 1576 -61
rect 1590 -64 1592 -61
rect 1497 -85 1499 -82
rect 1512 -85 1514 -82
rect 1528 -85 1530 -82
rect 1559 -85 1561 -82
rect 1590 -85 1592 -82
rect 1497 -125 1499 -95
rect 1512 -109 1514 -95
rect 1528 -125 1530 -95
rect 1543 -125 1545 -113
rect 1559 -125 1561 -95
rect 1574 -125 1576 -104
rect 1590 -125 1592 -95
rect 1497 -138 1499 -135
rect 1528 -138 1530 -135
rect 1543 -138 1545 -135
rect 1559 -138 1561 -135
rect 1574 -138 1576 -135
rect 1590 -138 1592 -135
rect 1274 -144 1279 -142
rect 1282 -144 1292 -142
rect 1296 -144 1309 -142
rect 1277 -145 1279 -144
rect 1290 -145 1292 -144
rect 1307 -145 1309 -144
rect 11 -162 13 -159
rect 26 -162 28 -159
rect 42 -162 44 -159
rect 73 -162 75 -159
rect 104 -162 106 -159
rect 1236 -158 1238 -155
rect 1260 -158 1262 -155
rect 1277 -158 1279 -155
rect 1290 -158 1292 -155
rect 1307 -158 1309 -155
rect 729 -161 731 -158
rect 743 -161 745 -158
rect 767 -161 769 -158
rect 791 -161 793 -158
rect 805 -161 807 -158
rect 829 -161 831 -158
rect 853 -161 855 -158
rect 867 -161 869 -158
rect 891 -161 893 -158
rect 1497 -159 1499 -156
rect 1512 -159 1514 -156
rect 1528 -159 1530 -156
rect 1559 -159 1561 -156
rect 1590 -159 1592 -156
rect 499 -168 501 -165
rect 513 -168 515 -165
rect 537 -168 539 -165
rect 561 -168 563 -165
rect 575 -168 577 -165
rect 599 -168 601 -165
rect 254 -171 256 -168
rect 268 -171 270 -168
rect 292 -171 294 -168
rect 11 -202 13 -172
rect 26 -186 28 -172
rect 42 -202 44 -172
rect 57 -202 59 -190
rect 73 -202 75 -172
rect 88 -202 90 -181
rect 104 -202 106 -172
rect 1236 -177 1238 -174
rect 1260 -177 1262 -174
rect 1274 -177 1276 -174
rect 1282 -177 1284 -174
rect 1296 -177 1298 -174
rect 11 -215 13 -212
rect 42 -215 44 -212
rect 57 -215 59 -212
rect 73 -215 75 -212
rect 88 -215 90 -212
rect 104 -215 106 -212
rect 254 -213 256 -191
rect 268 -213 270 -191
rect 292 -213 294 -191
rect 499 -198 501 -195
rect 513 -198 515 -195
rect 537 -198 539 -195
rect 1236 -212 1238 -197
rect 254 -226 256 -223
rect 268 -226 270 -223
rect 292 -226 294 -223
rect 11 -236 13 -233
rect 26 -236 28 -233
rect 42 -236 44 -233
rect 73 -236 75 -233
rect 104 -236 106 -233
rect 499 -240 501 -218
rect 513 -240 515 -218
rect 537 -240 539 -218
rect 1236 -225 1238 -222
rect 264 -245 266 -242
rect 288 -245 290 -242
rect 302 -245 304 -242
rect 310 -245 312 -242
rect 324 -245 326 -242
rect 11 -276 13 -246
rect 26 -260 28 -246
rect 42 -276 44 -246
rect 57 -276 59 -264
rect 73 -276 75 -246
rect 88 -276 90 -255
rect 104 -276 106 -246
rect 499 -253 501 -250
rect 513 -253 515 -250
rect 537 -253 539 -250
rect 1236 -260 1238 -257
rect 264 -280 266 -265
rect 11 -289 13 -286
rect 42 -289 44 -286
rect 57 -289 59 -286
rect 73 -289 75 -286
rect 88 -289 90 -286
rect 104 -289 106 -286
rect 264 -293 266 -290
rect 11 -310 13 -307
rect 26 -310 28 -307
rect 42 -310 44 -307
rect 73 -310 75 -307
rect 104 -310 106 -307
rect 11 -350 13 -320
rect 26 -334 28 -320
rect 42 -350 44 -320
rect 57 -350 59 -338
rect 73 -350 75 -320
rect 88 -350 90 -329
rect 104 -350 106 -320
rect 264 -328 266 -325
rect 11 -363 13 -360
rect 42 -363 44 -360
rect 57 -363 59 -360
rect 73 -363 75 -360
rect 88 -363 90 -360
rect 104 -363 106 -360
rect 264 -363 266 -348
rect 288 -363 290 -265
rect 302 -336 304 -265
rect 297 -338 304 -336
rect 297 -351 299 -338
rect 297 -353 304 -351
rect 302 -360 304 -353
rect 310 -360 312 -265
rect 324 -360 326 -265
rect 1236 -295 1238 -280
rect 1260 -295 1262 -197
rect 1274 -268 1276 -197
rect 1269 -270 1276 -268
rect 1269 -283 1271 -270
rect 1269 -285 1276 -283
rect 1274 -292 1276 -285
rect 1282 -292 1284 -197
rect 1296 -292 1298 -197
rect 1497 -199 1499 -169
rect 1512 -183 1514 -169
rect 1528 -199 1530 -169
rect 1543 -199 1545 -187
rect 1559 -199 1561 -169
rect 1574 -199 1576 -178
rect 1590 -199 1592 -169
rect 1497 -212 1499 -209
rect 1528 -212 1530 -209
rect 1543 -212 1545 -209
rect 1559 -212 1561 -209
rect 1574 -212 1576 -209
rect 1590 -212 1592 -209
rect 1497 -233 1499 -230
rect 1512 -233 1514 -230
rect 1528 -233 1530 -230
rect 1559 -233 1561 -230
rect 1590 -233 1592 -230
rect 1497 -273 1499 -243
rect 1512 -257 1514 -243
rect 1528 -273 1530 -243
rect 1543 -273 1545 -261
rect 1559 -273 1561 -243
rect 1574 -273 1576 -252
rect 1590 -273 1592 -243
rect 1497 -286 1499 -283
rect 1528 -286 1530 -283
rect 1543 -286 1545 -283
rect 1559 -286 1561 -283
rect 1574 -286 1576 -283
rect 1590 -286 1592 -283
rect 1274 -294 1279 -292
rect 1282 -294 1292 -292
rect 1296 -294 1309 -292
rect 1277 -295 1279 -294
rect 1290 -295 1292 -294
rect 1307 -295 1309 -294
rect 499 -310 501 -307
rect 513 -310 515 -307
rect 537 -310 539 -307
rect 561 -310 563 -307
rect 575 -310 577 -307
rect 599 -310 601 -307
rect 623 -310 625 -307
rect 637 -310 639 -307
rect 661 -310 663 -307
rect 685 -310 687 -307
rect 699 -310 701 -307
rect 723 -310 725 -307
rect 1236 -308 1238 -305
rect 1260 -308 1262 -305
rect 1277 -308 1279 -305
rect 1290 -308 1292 -305
rect 1307 -308 1309 -305
rect 1497 -307 1499 -304
rect 1512 -307 1514 -304
rect 1528 -307 1530 -304
rect 1559 -307 1561 -304
rect 1590 -307 1592 -304
rect 1236 -327 1238 -324
rect 1260 -327 1262 -324
rect 1274 -327 1276 -324
rect 1282 -327 1284 -324
rect 1296 -327 1298 -324
rect 499 -352 501 -330
rect 513 -352 515 -330
rect 537 -352 539 -330
rect 561 -352 563 -330
rect 575 -352 577 -330
rect 599 -352 601 -330
rect 623 -352 625 -330
rect 637 -352 639 -330
rect 661 -352 663 -330
rect 685 -352 687 -330
rect 699 -352 701 -330
rect 723 -352 725 -330
rect 1497 -347 1499 -317
rect 1512 -331 1514 -317
rect 1528 -347 1530 -317
rect 1543 -347 1545 -335
rect 1559 -347 1561 -317
rect 1574 -347 1576 -326
rect 1590 -347 1592 -317
rect 302 -362 307 -360
rect 310 -362 320 -360
rect 324 -362 337 -360
rect 1236 -362 1238 -347
rect 305 -363 307 -362
rect 318 -363 320 -362
rect 335 -363 337 -362
rect 499 -365 501 -362
rect 513 -365 515 -362
rect 537 -365 539 -362
rect 561 -365 563 -362
rect 575 -365 577 -362
rect 599 -365 601 -362
rect 623 -365 625 -362
rect 637 -365 639 -362
rect 661 -365 663 -362
rect 685 -365 687 -362
rect 699 -365 701 -362
rect 723 -365 725 -362
rect 264 -376 266 -373
rect 288 -376 290 -373
rect 305 -376 307 -373
rect 318 -376 320 -373
rect 335 -376 337 -373
rect 1236 -375 1238 -372
rect 11 -384 13 -381
rect 26 -384 28 -381
rect 42 -384 44 -381
rect 73 -384 75 -381
rect 104 -384 106 -381
rect 11 -424 13 -394
rect 26 -408 28 -394
rect 42 -424 44 -394
rect 57 -424 59 -412
rect 73 -424 75 -394
rect 88 -424 90 -403
rect 104 -424 106 -394
rect 254 -395 256 -392
rect 268 -395 270 -392
rect 292 -395 294 -392
rect 499 -410 501 -407
rect 513 -410 515 -407
rect 537 -410 539 -407
rect 561 -410 563 -407
rect 575 -410 577 -407
rect 599 -410 601 -407
rect 623 -410 625 -407
rect 637 -410 639 -407
rect 661 -410 663 -407
rect 1236 -410 1238 -407
rect 11 -437 13 -434
rect 42 -437 44 -434
rect 57 -437 59 -434
rect 73 -437 75 -434
rect 88 -437 90 -434
rect 104 -437 106 -434
rect 254 -437 256 -415
rect 268 -437 270 -415
rect 292 -437 294 -415
rect 254 -450 256 -447
rect 268 -450 270 -447
rect 292 -450 294 -447
rect 499 -452 501 -430
rect 513 -452 515 -430
rect 537 -452 539 -430
rect 561 -452 563 -430
rect 575 -452 577 -430
rect 599 -452 601 -430
rect 623 -452 625 -430
rect 637 -452 639 -430
rect 661 -452 663 -430
rect 1236 -445 1238 -430
rect 1260 -445 1262 -347
rect 1274 -418 1276 -347
rect 1269 -420 1276 -418
rect 1269 -433 1271 -420
rect 1269 -435 1276 -433
rect 1274 -442 1276 -435
rect 1282 -442 1284 -347
rect 1296 -442 1298 -347
rect 1497 -360 1499 -357
rect 1528 -360 1530 -357
rect 1543 -360 1545 -357
rect 1559 -360 1561 -357
rect 1574 -360 1576 -357
rect 1590 -360 1592 -357
rect 1274 -444 1279 -442
rect 1282 -444 1292 -442
rect 1296 -444 1309 -442
rect 1277 -445 1279 -444
rect 1290 -445 1292 -444
rect 1307 -445 1309 -444
rect 11 -458 13 -455
rect 26 -458 28 -455
rect 42 -458 44 -455
rect 73 -458 75 -455
rect 104 -458 106 -455
rect 1236 -458 1238 -455
rect 1260 -458 1262 -455
rect 1277 -458 1279 -455
rect 1290 -458 1292 -455
rect 1307 -458 1309 -455
rect 499 -465 501 -462
rect 513 -465 515 -462
rect 537 -465 539 -462
rect 561 -465 563 -462
rect 575 -465 577 -462
rect 599 -465 601 -462
rect 623 -465 625 -462
rect 637 -465 639 -462
rect 661 -465 663 -462
rect 11 -498 13 -468
rect 26 -482 28 -468
rect 42 -498 44 -468
rect 57 -498 59 -486
rect 73 -498 75 -468
rect 88 -498 90 -477
rect 104 -498 106 -468
rect 264 -469 266 -466
rect 288 -469 290 -466
rect 302 -469 304 -466
rect 310 -469 312 -466
rect 324 -469 326 -466
rect 264 -504 266 -489
rect 11 -511 13 -508
rect 42 -511 44 -508
rect 57 -511 59 -508
rect 73 -511 75 -508
rect 88 -511 90 -508
rect 104 -511 106 -508
rect 264 -517 266 -514
rect 264 -552 266 -549
rect 264 -587 266 -572
rect 288 -587 290 -489
rect 302 -560 304 -489
rect 297 -562 304 -560
rect 297 -575 299 -562
rect 297 -577 304 -575
rect 302 -584 304 -577
rect 310 -584 312 -489
rect 324 -584 326 -489
rect 807 -492 809 -489
rect 821 -492 823 -489
rect 845 -492 847 -489
rect 869 -492 871 -489
rect 883 -492 885 -489
rect 907 -492 909 -489
rect 931 -492 933 -489
rect 945 -492 947 -489
rect 969 -492 971 -489
rect 993 -492 995 -489
rect 1007 -492 1009 -489
rect 1031 -492 1033 -489
rect 499 -510 501 -507
rect 513 -510 515 -507
rect 537 -510 539 -507
rect 561 -510 563 -507
rect 575 -510 577 -507
rect 599 -510 601 -507
rect 499 -552 501 -530
rect 513 -552 515 -530
rect 537 -552 539 -530
rect 561 -552 563 -530
rect 575 -552 577 -530
rect 599 -552 601 -530
rect 807 -540 809 -512
rect 821 -540 823 -512
rect 845 -540 847 -512
rect 869 -540 871 -512
rect 883 -540 885 -512
rect 907 -540 909 -512
rect 931 -540 933 -512
rect 945 -540 947 -512
rect 969 -540 971 -512
rect 993 -540 995 -512
rect 1007 -540 1009 -512
rect 1031 -540 1033 -512
rect 807 -553 809 -550
rect 821 -553 823 -550
rect 845 -553 847 -550
rect 869 -553 871 -550
rect 883 -553 885 -550
rect 907 -553 909 -550
rect 931 -553 933 -550
rect 945 -553 947 -550
rect 969 -553 971 -550
rect 993 -553 995 -550
rect 1007 -553 1009 -550
rect 1031 -553 1033 -550
rect 499 -565 501 -562
rect 513 -565 515 -562
rect 537 -565 539 -562
rect 561 -565 563 -562
rect 575 -565 577 -562
rect 599 -565 601 -562
rect 302 -586 307 -584
rect 310 -586 320 -584
rect 324 -586 337 -584
rect 305 -587 307 -586
rect 318 -587 320 -586
rect 335 -587 337 -586
rect 264 -600 266 -597
rect 288 -600 290 -597
rect 305 -600 307 -597
rect 318 -600 320 -597
rect 335 -600 337 -597
rect 499 -610 501 -607
rect 513 -610 515 -607
rect 537 -610 539 -607
rect 254 -619 256 -616
rect 268 -619 270 -616
rect 292 -619 294 -616
rect 254 -661 256 -639
rect 268 -661 270 -639
rect 292 -661 294 -639
rect 499 -652 501 -630
rect 513 -652 515 -630
rect 537 -652 539 -630
rect 499 -665 501 -662
rect 513 -665 515 -662
rect 537 -665 539 -662
rect 254 -674 256 -671
rect 268 -674 270 -671
rect 292 -674 294 -671
<< polycontact >>
rect 495 216 499 220
rect 509 209 513 213
rect 533 216 537 220
rect 557 216 561 220
rect 571 209 575 213
rect 595 216 599 220
rect 260 172 264 176
rect 284 172 288 176
rect 260 89 264 93
rect 298 143 302 147
rect 495 127 499 131
rect 509 120 513 124
rect 533 127 537 131
rect 557 127 561 131
rect 571 120 575 124
rect 595 127 599 131
rect 1232 92 1236 96
rect 638 81 642 85
rect 652 74 656 78
rect 676 81 680 85
rect 700 81 704 85
rect 714 74 718 78
rect 738 81 742 85
rect 1256 92 1260 96
rect 6 28 11 33
rect 69 35 73 39
rect 53 28 57 32
rect 99 30 104 35
rect 495 44 499 48
rect 509 37 513 41
rect 533 44 537 48
rect 250 22 254 26
rect 264 15 268 19
rect 288 22 292 26
rect 1232 9 1236 13
rect 1270 63 1274 67
rect 6 -46 11 -41
rect 69 -39 73 -35
rect 53 -46 57 -42
rect 99 -44 104 -39
rect 260 -52 264 -48
rect 284 -52 288 -48
rect 6 -120 11 -115
rect 69 -113 73 -109
rect 53 -120 57 -116
rect 99 -118 104 -113
rect 260 -135 264 -131
rect 298 -81 302 -77
rect 495 -47 499 -43
rect 509 -54 513 -50
rect 533 -47 537 -43
rect 557 -47 561 -43
rect 571 -54 575 -50
rect 595 -47 599 -43
rect 619 -47 623 -43
rect 633 -54 637 -50
rect 657 -47 661 -43
rect 1492 -43 1497 -38
rect 1232 -58 1236 -54
rect 1256 -58 1260 -54
rect 725 -131 729 -127
rect 495 -144 499 -140
rect 509 -151 513 -147
rect 533 -144 537 -140
rect 557 -144 561 -140
rect 571 -151 575 -147
rect 595 -144 599 -140
rect 739 -138 743 -134
rect 763 -131 767 -127
rect 787 -131 791 -127
rect 801 -138 805 -134
rect 825 -131 829 -127
rect 849 -131 853 -127
rect 863 -138 867 -134
rect 887 -131 891 -127
rect 1232 -141 1236 -137
rect 1270 -87 1274 -83
rect 1555 -36 1559 -32
rect 1539 -43 1543 -39
rect 1585 -41 1590 -36
rect 1492 -117 1497 -112
rect 1555 -110 1559 -106
rect 1539 -117 1543 -113
rect 1585 -115 1590 -110
rect 6 -194 11 -189
rect 69 -187 73 -183
rect 53 -194 57 -190
rect 99 -192 104 -187
rect 250 -202 254 -198
rect 264 -209 268 -205
rect 288 -202 292 -198
rect 1492 -191 1497 -186
rect 1232 -208 1236 -204
rect 1256 -208 1260 -204
rect 495 -229 499 -225
rect 509 -236 513 -232
rect 533 -229 537 -225
rect 6 -268 11 -263
rect 69 -261 73 -257
rect 53 -268 57 -264
rect 99 -266 104 -261
rect 260 -276 264 -272
rect 284 -276 288 -272
rect 6 -342 11 -337
rect 69 -335 73 -331
rect 53 -342 57 -338
rect 99 -340 104 -335
rect 260 -359 264 -355
rect 298 -305 302 -301
rect 1232 -291 1236 -287
rect 1270 -237 1274 -233
rect 1555 -184 1559 -180
rect 1539 -191 1543 -187
rect 1585 -189 1590 -184
rect 1492 -265 1497 -260
rect 1555 -258 1559 -254
rect 1539 -265 1543 -261
rect 1585 -263 1590 -258
rect 495 -341 499 -337
rect 509 -348 513 -344
rect 533 -341 537 -337
rect 557 -341 561 -337
rect 571 -348 575 -344
rect 595 -341 599 -337
rect 619 -341 623 -337
rect 633 -348 637 -344
rect 657 -341 661 -337
rect 681 -341 685 -337
rect 695 -348 699 -344
rect 719 -341 723 -337
rect 1492 -339 1497 -334
rect 1555 -332 1559 -328
rect 1539 -339 1543 -335
rect 1585 -337 1590 -332
rect 1232 -358 1236 -354
rect 1256 -358 1260 -354
rect 6 -416 11 -411
rect 69 -409 73 -405
rect 53 -416 57 -412
rect 99 -414 104 -409
rect 250 -426 254 -422
rect 264 -433 268 -429
rect 288 -426 292 -422
rect 495 -441 499 -437
rect 509 -448 513 -444
rect 533 -441 537 -437
rect 557 -441 561 -437
rect 571 -448 575 -444
rect 595 -441 599 -437
rect 619 -441 623 -437
rect 633 -448 637 -444
rect 657 -441 661 -437
rect 1232 -441 1236 -437
rect 1270 -387 1274 -383
rect 6 -490 11 -485
rect 69 -483 73 -479
rect 53 -490 57 -486
rect 99 -488 104 -483
rect 260 -500 264 -496
rect 284 -500 288 -496
rect 260 -583 264 -579
rect 298 -529 302 -525
rect 803 -523 807 -519
rect 495 -541 499 -537
rect 509 -548 513 -544
rect 533 -541 537 -537
rect 557 -541 561 -537
rect 571 -548 575 -544
rect 595 -541 599 -537
rect 817 -530 821 -526
rect 841 -523 845 -519
rect 865 -523 869 -519
rect 879 -530 883 -526
rect 903 -523 907 -519
rect 927 -523 931 -519
rect 941 -530 945 -526
rect 965 -523 969 -519
rect 989 -523 993 -519
rect 1003 -530 1007 -526
rect 1027 -523 1031 -519
rect 250 -650 254 -646
rect 264 -657 268 -653
rect 288 -650 292 -646
rect 495 -641 499 -637
rect 509 -648 513 -644
rect 533 -641 537 -637
<< metal1 >>
rect 405 305 1205 310
rect 405 213 410 305
rect 473 279 1165 283
rect 473 220 477 279
rect 494 255 607 257
rect 494 251 536 255
rect 540 251 598 255
rect 602 251 607 255
rect 494 247 498 251
rect 516 247 520 251
rect 532 247 536 251
rect 556 247 560 251
rect 594 247 598 251
rect 505 220 509 227
rect 540 220 544 227
rect 578 220 582 227
rect 602 220 606 227
rect 473 216 495 220
rect 505 216 533 220
rect 540 216 557 220
rect 578 216 595 220
rect 602 216 1117 220
rect 253 211 277 213
rect 253 207 263 211
rect 267 207 277 211
rect 282 207 326 213
rect 259 203 263 207
rect 283 203 287 207
rect 327 203 331 207
rect 405 208 463 213
rect 267 176 271 183
rect 239 172 260 176
rect 267 172 284 176
rect 239 146 243 172
rect 267 168 271 172
rect 259 154 263 158
rect 251 149 263 154
rect 266 150 296 154
rect 266 146 270 150
rect 145 142 270 146
rect 273 143 298 147
rect 145 141 234 142
rect 0 68 103 70
rect 0 64 54 68
rect 58 64 103 68
rect 6 60 10 64
rect 37 60 41 64
rect 68 60 72 64
rect 99 60 103 64
rect -23 36 3 41
rect -23 -33 -18 36
rect 0 28 6 33
rect 29 32 33 50
rect 45 39 49 50
rect 76 48 80 50
rect 76 44 95 48
rect 45 35 69 39
rect 91 35 95 44
rect 107 35 111 50
rect 145 35 150 141
rect 14 28 53 32
rect 14 20 18 28
rect 60 20 64 35
rect 91 30 99 35
rect 107 30 150 35
rect 174 89 220 94
rect 91 20 95 30
rect 107 20 111 30
rect 6 6 10 10
rect 37 6 41 10
rect 68 6 72 10
rect 99 6 103 10
rect 0 4 103 6
rect 0 0 52 4
rect 56 0 103 4
rect 0 -6 103 -4
rect 0 -10 54 -6
rect 58 -10 103 -6
rect 6 -14 10 -10
rect 37 -14 41 -10
rect 68 -14 72 -10
rect 99 -14 103 -10
rect -23 -38 3 -33
rect -23 -107 -18 -38
rect 0 -46 6 -41
rect 29 -42 33 -24
rect 45 -35 49 -24
rect 76 -26 80 -24
rect 76 -30 95 -26
rect 45 -39 69 -35
rect 91 -39 95 -30
rect 107 -39 111 -24
rect 174 -39 179 89
rect 230 19 234 141
rect 273 138 277 143
rect 305 140 309 183
rect 405 140 409 208
rect 246 134 277 138
rect 283 136 409 140
rect 246 93 250 134
rect 253 128 272 130
rect 253 124 263 128
rect 267 124 272 128
rect 259 120 263 124
rect 267 93 271 100
rect 242 89 260 93
rect 239 26 243 89
rect 267 88 272 93
rect 267 85 271 88
rect 283 85 287 136
rect 291 88 325 92
rect 291 85 295 88
rect 321 85 325 88
rect 338 85 342 136
rect 473 131 477 216
rect 492 209 509 213
rect 516 205 520 216
rect 540 205 544 216
rect 553 209 571 213
rect 578 206 582 216
rect 556 202 582 206
rect 556 199 560 202
rect 578 199 582 202
rect 602 199 606 216
rect 494 191 498 195
rect 532 191 536 195
rect 494 187 504 191
rect 509 187 536 191
rect 540 187 548 191
rect 544 185 548 187
rect 567 185 571 189
rect 594 185 598 189
rect 544 181 598 185
rect 602 181 629 185
rect 488 172 548 177
rect 494 166 607 168
rect 494 162 536 166
rect 540 162 598 166
rect 602 162 607 166
rect 494 158 498 162
rect 516 158 520 162
rect 532 158 536 162
rect 556 158 560 162
rect 578 158 582 162
rect 594 158 598 162
rect 505 131 509 138
rect 540 131 544 138
rect 567 131 571 138
rect 602 131 606 138
rect 473 127 495 131
rect 505 127 533 131
rect 540 127 557 131
rect 567 127 595 131
rect 602 127 623 131
rect 259 72 263 75
rect 251 67 263 72
rect 310 71 314 75
rect 267 67 314 71
rect 249 61 300 63
rect 249 57 291 61
rect 295 57 300 61
rect 249 53 253 57
rect 271 53 275 57
rect 287 53 291 57
rect 260 26 264 33
rect 295 26 299 33
rect 239 22 250 26
rect 260 22 288 26
rect 295 22 351 26
rect 230 15 264 19
rect 271 11 275 22
rect 295 11 299 22
rect 249 -2 253 1
rect 251 -3 253 -2
rect 287 -3 291 1
rect 251 -7 291 -3
rect 253 -13 277 -11
rect 253 -17 263 -13
rect 267 -17 277 -13
rect 282 -17 326 -11
rect 14 -46 53 -42
rect 14 -54 18 -46
rect 60 -54 64 -39
rect 91 -44 99 -39
rect 107 -44 179 -39
rect 259 -21 263 -17
rect 283 -21 287 -17
rect 327 -21 331 -17
rect 91 -54 95 -44
rect 107 -54 111 -44
rect 267 -48 271 -41
rect 239 -52 260 -48
rect 267 -52 284 -48
rect 6 -68 10 -64
rect 37 -68 41 -64
rect 68 -68 72 -64
rect 99 -68 103 -64
rect 0 -70 103 -68
rect 0 -74 52 -70
rect 56 -74 103 -70
rect 239 -78 243 -52
rect 267 -56 271 -52
rect 259 -70 263 -66
rect 251 -75 263 -70
rect 266 -74 296 -70
rect 266 -78 270 -74
rect 0 -80 103 -78
rect 0 -84 54 -80
rect 58 -84 103 -80
rect 6 -88 10 -84
rect 37 -88 41 -84
rect 68 -88 72 -84
rect 99 -88 103 -84
rect 166 -82 270 -78
rect 273 -81 298 -77
rect 166 -83 234 -82
rect -23 -112 3 -107
rect -23 -181 -18 -112
rect 0 -120 6 -115
rect 29 -116 33 -98
rect 45 -109 49 -98
rect 76 -100 80 -98
rect 76 -104 95 -100
rect 45 -113 69 -109
rect 91 -113 95 -104
rect 107 -113 111 -98
rect 166 -113 171 -83
rect 14 -120 53 -116
rect 14 -128 18 -120
rect 60 -128 64 -113
rect 91 -118 99 -113
rect 107 -118 171 -113
rect 91 -128 95 -118
rect 107 -128 111 -118
rect 183 -135 220 -130
rect 6 -142 10 -138
rect 37 -142 41 -138
rect 68 -142 72 -138
rect 99 -142 103 -138
rect 0 -144 103 -142
rect 0 -148 52 -144
rect 56 -148 103 -144
rect 0 -154 103 -152
rect 0 -158 54 -154
rect 58 -158 103 -154
rect 6 -162 10 -158
rect 37 -162 41 -158
rect 68 -162 72 -158
rect 99 -162 103 -158
rect -23 -186 3 -181
rect -23 -255 -18 -186
rect 0 -194 6 -189
rect 29 -190 33 -172
rect 45 -183 49 -172
rect 76 -174 80 -172
rect 76 -178 95 -174
rect 45 -187 69 -183
rect 91 -187 95 -178
rect 107 -187 111 -172
rect 183 -187 188 -135
rect 14 -194 53 -190
rect 14 -202 18 -194
rect 60 -202 64 -187
rect 91 -192 99 -187
rect 107 -192 188 -187
rect 91 -202 95 -192
rect 107 -202 111 -192
rect 230 -205 234 -83
rect 273 -86 277 -81
rect 305 -84 309 -41
rect 473 -43 477 127
rect 488 123 509 124
rect 491 120 509 123
rect 516 116 520 127
rect 540 116 544 127
rect 554 120 571 124
rect 578 116 582 127
rect 602 116 606 127
rect 494 102 498 106
rect 494 98 504 102
rect 532 102 536 106
rect 556 102 560 106
rect 594 102 598 106
rect 509 98 536 102
rect 540 98 598 102
rect 602 98 612 102
rect 485 89 549 94
rect 485 48 490 89
rect 619 85 623 127
rect 631 116 641 122
rect 647 120 755 122
rect 647 116 679 120
rect 683 116 741 120
rect 745 116 755 120
rect 637 112 641 116
rect 675 112 679 116
rect 699 112 703 116
rect 737 112 741 116
rect 659 85 663 92
rect 683 85 687 92
rect 721 85 725 92
rect 745 85 749 92
rect 494 83 544 85
rect 494 79 536 83
rect 540 79 544 83
rect 619 81 638 85
rect 659 81 676 85
rect 683 81 700 85
rect 721 81 738 85
rect 745 81 1073 85
rect 494 75 498 79
rect 516 75 520 79
rect 532 75 536 79
rect 505 48 509 55
rect 540 48 544 55
rect 619 74 652 78
rect 619 48 623 74
rect 659 71 663 81
rect 637 67 663 71
rect 637 64 641 67
rect 659 64 663 67
rect 683 64 687 81
rect 696 74 714 78
rect 721 71 725 81
rect 699 67 725 71
rect 699 64 703 67
rect 721 64 725 67
rect 745 64 749 81
rect 485 44 495 48
rect 505 44 533 48
rect 540 44 623 48
rect 648 50 652 54
rect 675 50 679 54
rect 710 50 714 54
rect 737 50 741 54
rect 648 46 679 50
rect 683 46 741 50
rect 745 46 750 50
rect 488 37 509 41
rect 516 33 520 44
rect 540 33 544 44
rect 659 37 691 42
rect 494 19 498 23
rect 494 15 504 19
rect 532 19 536 23
rect 509 15 536 19
rect 494 -8 616 -6
rect 494 -12 536 -8
rect 540 -12 598 -8
rect 602 -12 616 -8
rect 622 -8 674 -6
rect 622 -12 660 -8
rect 664 -12 674 -8
rect 494 -16 498 -12
rect 516 -16 520 -12
rect 532 -16 536 -12
rect 556 -16 560 -12
rect 578 -16 582 -12
rect 594 -16 598 -12
rect 618 -16 622 -12
rect 640 -16 644 -12
rect 656 -16 660 -12
rect 505 -43 509 -36
rect 540 -43 544 -36
rect 567 -43 571 -36
rect 602 -43 606 -36
rect 629 -43 633 -36
rect 664 -43 668 -36
rect 473 -47 495 -43
rect 505 -47 533 -43
rect 540 -47 557 -43
rect 567 -47 595 -43
rect 602 -47 619 -43
rect 629 -47 657 -43
rect 664 -47 697 -43
rect 246 -90 277 -86
rect 283 -88 351 -84
rect 246 -131 250 -90
rect 253 -96 272 -94
rect 253 -100 263 -96
rect 267 -100 272 -96
rect 259 -104 263 -100
rect 267 -131 271 -124
rect 242 -135 260 -131
rect 239 -198 243 -135
rect 267 -136 272 -131
rect 267 -139 271 -136
rect 283 -139 287 -88
rect 291 -136 325 -132
rect 291 -139 295 -136
rect 321 -139 325 -136
rect 338 -139 342 -88
rect 259 -152 263 -149
rect 251 -157 263 -152
rect 310 -153 314 -149
rect 267 -157 314 -153
rect 249 -163 300 -161
rect 249 -167 291 -163
rect 295 -167 300 -163
rect 249 -171 253 -167
rect 271 -171 275 -167
rect 287 -171 291 -167
rect 260 -198 264 -191
rect 295 -198 299 -191
rect 239 -202 250 -198
rect 260 -202 288 -198
rect 295 -202 351 -198
rect 230 -209 264 -205
rect 6 -216 10 -212
rect 37 -216 41 -212
rect 68 -216 72 -212
rect 99 -216 103 -212
rect 271 -213 275 -202
rect 295 -213 299 -202
rect 0 -218 103 -216
rect 0 -222 52 -218
rect 56 -222 103 -218
rect 249 -226 253 -223
rect 0 -228 103 -226
rect 0 -232 54 -228
rect 58 -232 103 -228
rect 251 -227 253 -226
rect 287 -227 291 -223
rect 251 -231 291 -227
rect 6 -236 10 -232
rect 37 -236 41 -232
rect 68 -236 72 -232
rect 99 -236 103 -232
rect 253 -237 277 -235
rect 253 -241 263 -237
rect 267 -241 277 -237
rect 282 -241 326 -235
rect -23 -260 3 -255
rect -23 -329 -18 -260
rect 0 -268 6 -263
rect 29 -264 33 -246
rect 45 -257 49 -246
rect 76 -248 80 -246
rect 76 -252 95 -248
rect 45 -261 69 -257
rect 91 -261 95 -252
rect 107 -261 111 -246
rect 259 -245 263 -241
rect 283 -245 287 -241
rect 327 -245 331 -241
rect 14 -268 53 -264
rect 14 -276 18 -268
rect 60 -276 64 -261
rect 91 -266 99 -261
rect 107 -266 193 -261
rect 91 -276 95 -266
rect 107 -276 111 -266
rect 6 -290 10 -286
rect 37 -290 41 -286
rect 68 -290 72 -286
rect 99 -290 103 -286
rect 0 -292 103 -290
rect 0 -296 52 -292
rect 56 -296 103 -292
rect 0 -302 103 -300
rect 0 -306 54 -302
rect 58 -306 103 -302
rect 6 -310 10 -306
rect 37 -310 41 -306
rect 68 -310 72 -306
rect 99 -310 103 -306
rect 188 -302 193 -266
rect 267 -272 271 -265
rect 239 -276 260 -272
rect 267 -276 284 -272
rect 239 -302 243 -276
rect 267 -280 271 -276
rect 259 -294 263 -290
rect 251 -299 263 -294
rect 266 -298 296 -294
rect 266 -302 270 -298
rect 188 -306 270 -302
rect 273 -305 298 -301
rect 188 -307 234 -306
rect -23 -334 3 -329
rect -23 -403 -18 -334
rect 0 -342 6 -337
rect 29 -338 33 -320
rect 45 -331 49 -320
rect 76 -322 80 -320
rect 76 -326 95 -322
rect 45 -335 69 -331
rect 91 -335 95 -326
rect 107 -335 111 -320
rect 14 -342 53 -338
rect 14 -350 18 -342
rect 60 -350 64 -335
rect 91 -340 99 -335
rect 107 -340 194 -335
rect 91 -350 95 -340
rect 107 -350 111 -340
rect 189 -354 194 -340
rect 189 -359 220 -354
rect 6 -364 10 -360
rect 37 -364 41 -360
rect 68 -364 72 -360
rect 99 -364 103 -360
rect 0 -366 103 -364
rect 0 -370 52 -366
rect 56 -370 103 -366
rect 0 -376 103 -374
rect 0 -380 54 -376
rect 58 -380 103 -376
rect 6 -384 10 -380
rect 37 -384 41 -380
rect 68 -384 72 -380
rect 99 -384 103 -380
rect -23 -408 3 -403
rect -23 -477 -18 -408
rect 0 -416 6 -411
rect 29 -412 33 -394
rect 45 -405 49 -394
rect 76 -396 80 -394
rect 76 -400 95 -396
rect 45 -409 69 -405
rect 91 -409 95 -400
rect 107 -409 111 -394
rect 14 -416 53 -412
rect 14 -424 18 -416
rect 60 -424 64 -409
rect 91 -414 99 -409
rect 107 -414 187 -409
rect 91 -424 95 -414
rect 107 -424 111 -414
rect 6 -438 10 -434
rect 37 -438 41 -434
rect 68 -438 72 -434
rect 99 -438 103 -434
rect 0 -440 103 -438
rect 0 -444 52 -440
rect 56 -444 103 -440
rect 0 -450 103 -448
rect 0 -454 54 -450
rect 58 -454 103 -450
rect 6 -458 10 -454
rect 37 -458 41 -454
rect 68 -458 72 -454
rect 99 -458 103 -454
rect -23 -482 3 -477
rect -23 -748 -18 -482
rect 0 -490 6 -485
rect 29 -486 33 -468
rect 45 -479 49 -468
rect 76 -470 80 -468
rect 76 -474 95 -470
rect 45 -483 69 -479
rect 91 -483 95 -474
rect 107 -483 111 -468
rect 14 -490 53 -486
rect 14 -498 18 -490
rect 60 -498 64 -483
rect 91 -488 99 -483
rect 107 -488 151 -483
rect 91 -498 95 -488
rect 107 -498 111 -488
rect 6 -512 10 -508
rect 37 -512 41 -508
rect 68 -512 72 -508
rect 99 -512 103 -508
rect 0 -514 103 -512
rect 0 -518 52 -514
rect 56 -518 103 -514
rect 146 -578 151 -488
rect 182 -526 187 -414
rect 230 -429 234 -307
rect 273 -310 277 -305
rect 305 -308 309 -265
rect 246 -314 277 -310
rect 283 -312 351 -308
rect 246 -355 250 -314
rect 253 -320 272 -318
rect 253 -324 263 -320
rect 267 -324 272 -320
rect 259 -328 263 -324
rect 267 -355 271 -348
rect 242 -359 260 -355
rect 239 -422 243 -359
rect 267 -360 272 -355
rect 267 -363 271 -360
rect 283 -363 287 -312
rect 291 -360 325 -356
rect 291 -363 295 -360
rect 321 -363 325 -360
rect 338 -363 342 -312
rect 473 -337 477 -47
rect 486 -51 509 -50
rect 490 -54 509 -51
rect 516 -58 520 -47
rect 540 -58 544 -47
rect 553 -54 571 -50
rect 578 -58 582 -47
rect 602 -58 606 -47
rect 616 -54 633 -50
rect 640 -58 644 -47
rect 664 -58 668 -47
rect 494 -72 498 -68
rect 494 -76 504 -72
rect 532 -72 536 -68
rect 556 -72 560 -68
rect 594 -72 598 -68
rect 618 -72 622 -68
rect 656 -72 660 -68
rect 509 -76 536 -72
rect 540 -76 598 -72
rect 602 -76 660 -72
rect 664 -76 674 -72
rect 481 -85 548 -80
rect 602 -85 611 -80
rect 481 -140 486 -85
rect 494 -105 607 -103
rect 494 -109 536 -105
rect 540 -109 598 -105
rect 602 -109 607 -105
rect 494 -113 498 -109
rect 516 -113 520 -109
rect 532 -113 536 -109
rect 556 -113 560 -109
rect 578 -113 582 -109
rect 594 -113 598 -109
rect 693 -127 697 -47
rect 718 -96 719 -90
rect 725 -92 904 -90
rect 725 -96 766 -92
rect 770 -96 828 -92
rect 832 -96 890 -92
rect 894 -96 904 -92
rect 724 -100 728 -96
rect 762 -100 766 -96
rect 786 -100 790 -96
rect 824 -100 828 -96
rect 848 -100 852 -96
rect 886 -100 890 -96
rect 746 -127 750 -120
rect 770 -127 774 -120
rect 808 -127 812 -120
rect 832 -127 836 -120
rect 870 -127 874 -120
rect 894 -127 898 -120
rect 693 -131 725 -127
rect 746 -131 763 -127
rect 770 -131 787 -127
rect 808 -131 825 -127
rect 832 -131 849 -127
rect 870 -131 887 -127
rect 894 -131 1023 -127
rect 505 -140 509 -133
rect 540 -140 544 -133
rect 567 -140 571 -133
rect 602 -140 606 -133
rect 693 -138 739 -134
rect 693 -140 697 -138
rect 481 -144 495 -140
rect 505 -144 533 -140
rect 540 -144 557 -140
rect 567 -144 595 -140
rect 602 -144 697 -140
rect 746 -141 750 -131
rect 488 -151 509 -147
rect 516 -155 520 -144
rect 540 -155 544 -144
rect 553 -151 571 -147
rect 578 -155 582 -144
rect 602 -155 606 -144
rect 724 -145 750 -141
rect 724 -148 728 -145
rect 746 -148 750 -145
rect 770 -148 774 -131
rect 783 -138 801 -134
rect 808 -141 812 -131
rect 786 -145 812 -141
rect 786 -148 790 -145
rect 808 -148 812 -145
rect 832 -148 836 -131
rect 845 -138 863 -134
rect 870 -141 874 -131
rect 848 -145 874 -141
rect 848 -148 852 -145
rect 870 -148 874 -145
rect 894 -148 898 -131
rect 735 -162 739 -158
rect 762 -162 766 -158
rect 797 -162 801 -158
rect 824 -162 828 -158
rect 859 -162 863 -158
rect 886 -162 890 -158
rect 494 -169 498 -165
rect 494 -173 504 -169
rect 532 -169 536 -165
rect 556 -169 560 -165
rect 594 -169 598 -165
rect 721 -166 766 -162
rect 770 -166 828 -162
rect 832 -166 890 -162
rect 894 -166 899 -162
rect 509 -173 536 -169
rect 540 -173 598 -169
rect 602 -173 612 -169
rect 727 -175 778 -170
rect 833 -175 840 -170
rect 540 -182 548 -177
rect 494 -190 545 -188
rect 494 -194 536 -190
rect 540 -194 545 -190
rect 494 -198 498 -194
rect 516 -198 520 -194
rect 532 -198 536 -194
rect 505 -225 509 -218
rect 540 -225 544 -218
rect 727 -225 731 -175
rect 488 -229 495 -225
rect 505 -229 533 -225
rect 540 -229 731 -225
rect 488 -236 509 -232
rect 516 -240 520 -229
rect 540 -240 544 -229
rect 494 -254 498 -250
rect 494 -258 504 -254
rect 532 -254 536 -250
rect 509 -258 536 -254
rect 540 -258 548 -254
rect 494 -302 681 -300
rect 494 -306 536 -302
rect 540 -306 598 -302
rect 602 -306 660 -302
rect 664 -306 681 -302
rect 687 -302 736 -300
rect 687 -306 722 -302
rect 726 -306 736 -302
rect 494 -310 498 -306
rect 516 -310 520 -306
rect 532 -310 536 -306
rect 556 -310 560 -306
rect 578 -310 582 -306
rect 594 -310 598 -306
rect 618 -310 622 -306
rect 640 -310 644 -306
rect 656 -310 660 -306
rect 680 -310 684 -306
rect 702 -310 706 -306
rect 718 -310 722 -306
rect 505 -337 509 -330
rect 540 -337 544 -330
rect 567 -337 571 -330
rect 602 -337 606 -330
rect 629 -337 633 -330
rect 664 -337 668 -330
rect 691 -337 695 -330
rect 726 -337 730 -330
rect 473 -341 495 -337
rect 505 -341 533 -337
rect 540 -341 557 -337
rect 567 -341 595 -337
rect 602 -341 619 -337
rect 629 -341 657 -337
rect 664 -341 681 -337
rect 691 -341 719 -337
rect 726 -341 752 -337
rect 491 -348 509 -344
rect 516 -352 520 -341
rect 540 -352 544 -341
rect 554 -348 571 -344
rect 578 -352 582 -341
rect 602 -352 606 -341
rect 615 -348 633 -344
rect 640 -352 644 -341
rect 664 -352 668 -341
rect 677 -348 695 -344
rect 702 -352 706 -341
rect 726 -352 730 -341
rect 494 -366 498 -362
rect 494 -370 504 -366
rect 532 -366 536 -362
rect 556 -366 560 -362
rect 594 -366 598 -362
rect 618 -366 622 -362
rect 656 -366 660 -362
rect 680 -366 684 -362
rect 718 -366 722 -362
rect 509 -370 536 -366
rect 540 -370 598 -366
rect 602 -370 660 -366
rect 664 -370 722 -366
rect 726 -370 736 -366
rect 259 -376 263 -373
rect 251 -381 263 -376
rect 310 -377 314 -373
rect 267 -381 314 -377
rect 544 -379 549 -374
rect 604 -379 610 -374
rect 666 -379 672 -374
rect 249 -387 300 -385
rect 249 -391 291 -387
rect 295 -391 300 -387
rect 249 -395 253 -391
rect 271 -395 275 -391
rect 287 -395 291 -391
rect 260 -422 264 -415
rect 295 -422 299 -415
rect 494 -402 669 -400
rect 494 -406 536 -402
rect 540 -406 598 -402
rect 602 -406 660 -402
rect 664 -406 669 -402
rect 494 -410 498 -406
rect 516 -410 520 -406
rect 239 -426 250 -422
rect 260 -426 288 -422
rect 295 -426 351 -422
rect 230 -433 264 -429
rect 271 -437 275 -426
rect 295 -437 299 -426
rect 532 -410 536 -406
rect 556 -410 560 -406
rect 578 -410 582 -406
rect 594 -410 598 -406
rect 618 -410 622 -406
rect 640 -410 644 -406
rect 656 -410 660 -406
rect 505 -437 509 -430
rect 540 -437 544 -430
rect 567 -437 571 -430
rect 602 -437 606 -430
rect 629 -437 633 -430
rect 664 -437 668 -430
rect 488 -441 495 -437
rect 505 -441 533 -437
rect 540 -441 557 -437
rect 567 -441 595 -437
rect 602 -441 619 -437
rect 629 -441 657 -437
rect 664 -441 721 -437
rect 249 -450 253 -447
rect 251 -451 253 -450
rect 287 -451 291 -447
rect 488 -448 509 -444
rect 251 -455 291 -451
rect 516 -452 520 -441
rect 540 -452 544 -441
rect 554 -448 571 -444
rect 578 -452 582 -441
rect 602 -452 606 -441
rect 615 -448 633 -444
rect 640 -452 644 -441
rect 664 -452 668 -441
rect 253 -461 277 -459
rect 253 -465 263 -461
rect 267 -465 277 -461
rect 282 -465 326 -459
rect 259 -469 263 -465
rect 283 -469 287 -465
rect 327 -469 331 -465
rect 494 -466 498 -462
rect 494 -470 504 -466
rect 532 -466 536 -462
rect 556 -466 560 -462
rect 594 -466 598 -462
rect 618 -466 622 -462
rect 656 -466 660 -462
rect 509 -470 536 -466
rect 540 -470 598 -466
rect 602 -470 660 -466
rect 664 -470 674 -466
rect 544 -479 549 -474
rect 604 -479 610 -474
rect 267 -496 271 -489
rect 239 -500 260 -496
rect 267 -500 284 -496
rect 239 -526 243 -500
rect 267 -504 271 -500
rect 259 -518 263 -514
rect 251 -523 263 -518
rect 266 -522 296 -518
rect 266 -526 270 -522
rect 182 -530 270 -526
rect 273 -529 298 -525
rect 182 -531 234 -530
rect 146 -583 220 -578
rect 230 -653 234 -531
rect 273 -534 277 -529
rect 305 -532 309 -489
rect 494 -502 607 -500
rect 494 -506 536 -502
rect 540 -506 598 -502
rect 602 -506 607 -502
rect 494 -510 498 -506
rect 516 -510 520 -506
rect 532 -510 536 -506
rect 556 -510 560 -506
rect 578 -510 582 -506
rect 594 -510 598 -506
rect 717 -526 721 -441
rect 748 -519 752 -341
rect 1019 -437 1023 -131
rect 1069 -287 1073 81
rect 1113 -137 1117 216
rect 1161 13 1165 279
rect 1200 96 1205 305
rect 1225 131 1249 133
rect 1225 127 1235 131
rect 1239 127 1249 131
rect 1254 127 1303 133
rect 1231 123 1235 127
rect 1255 123 1259 127
rect 1299 123 1303 127
rect 1239 96 1243 103
rect 1200 92 1232 96
rect 1239 92 1256 96
rect 1200 91 1216 92
rect 1211 66 1215 91
rect 1239 88 1243 92
rect 1231 74 1235 78
rect 1223 69 1235 74
rect 1238 70 1268 74
rect 1238 66 1242 70
rect 1211 62 1242 66
rect 1245 63 1270 67
rect 1245 58 1249 63
rect 1277 60 1281 103
rect 1218 54 1249 58
rect 1255 56 1447 60
rect 1218 13 1222 54
rect 1225 48 1244 50
rect 1225 44 1235 48
rect 1239 44 1244 48
rect 1231 40 1235 44
rect 1239 13 1243 20
rect 1161 9 1232 13
rect 1239 8 1244 13
rect 1239 5 1243 8
rect 1255 5 1259 56
rect 1263 8 1297 12
rect 1263 5 1267 8
rect 1293 5 1297 8
rect 1310 5 1314 56
rect 1231 -8 1235 -5
rect 1223 -13 1235 -8
rect 1282 -9 1286 -5
rect 1239 -13 1286 -9
rect 1225 -19 1249 -17
rect 1225 -23 1235 -19
rect 1239 -23 1249 -19
rect 1254 -23 1303 -17
rect 1231 -27 1235 -23
rect 1255 -27 1259 -23
rect 1299 -27 1303 -23
rect 1443 -38 1447 56
rect 1486 -3 1589 -1
rect 1486 -7 1540 -3
rect 1544 -7 1589 -3
rect 1492 -11 1496 -7
rect 1523 -11 1527 -7
rect 1554 -11 1558 -7
rect 1585 -11 1589 -7
rect 1443 -43 1492 -38
rect 1515 -39 1519 -21
rect 1531 -32 1535 -21
rect 1562 -23 1566 -21
rect 1562 -27 1581 -23
rect 1531 -36 1555 -32
rect 1577 -36 1581 -27
rect 1593 -36 1597 -21
rect 1500 -43 1539 -39
rect 1239 -54 1243 -47
rect 1211 -58 1232 -54
rect 1239 -58 1256 -54
rect 1211 -84 1215 -58
rect 1239 -62 1243 -58
rect 1231 -76 1235 -72
rect 1223 -81 1235 -76
rect 1238 -80 1268 -76
rect 1238 -84 1242 -80
rect 1211 -88 1242 -84
rect 1245 -87 1270 -83
rect 1245 -92 1249 -87
rect 1277 -90 1281 -47
rect 1500 -51 1504 -43
rect 1546 -51 1550 -36
rect 1577 -41 1585 -36
rect 1593 -41 1608 -36
rect 1577 -51 1581 -41
rect 1593 -51 1597 -41
rect 1492 -65 1496 -61
rect 1523 -65 1527 -61
rect 1554 -65 1558 -61
rect 1585 -65 1589 -61
rect 1486 -67 1589 -65
rect 1486 -71 1538 -67
rect 1542 -71 1589 -67
rect 1486 -77 1589 -75
rect 1486 -81 1540 -77
rect 1544 -81 1589 -77
rect 1492 -85 1496 -81
rect 1523 -85 1527 -81
rect 1554 -85 1558 -81
rect 1585 -85 1589 -81
rect 1218 -96 1249 -92
rect 1255 -94 1449 -90
rect 1218 -137 1222 -96
rect 1225 -102 1244 -100
rect 1225 -106 1235 -102
rect 1239 -106 1244 -102
rect 1231 -110 1235 -106
rect 1239 -137 1243 -130
rect 1113 -141 1232 -137
rect 1239 -142 1244 -137
rect 1239 -145 1243 -142
rect 1255 -145 1259 -94
rect 1263 -142 1297 -138
rect 1263 -145 1267 -142
rect 1293 -145 1297 -142
rect 1310 -145 1314 -94
rect 1445 -112 1449 -94
rect 1445 -117 1492 -112
rect 1515 -113 1519 -95
rect 1531 -106 1535 -95
rect 1562 -97 1566 -95
rect 1562 -101 1581 -97
rect 1531 -110 1555 -106
rect 1577 -110 1581 -101
rect 1593 -110 1597 -95
rect 1500 -117 1539 -113
rect 1500 -125 1504 -117
rect 1546 -125 1550 -110
rect 1577 -115 1585 -110
rect 1593 -115 1608 -110
rect 1577 -125 1581 -115
rect 1593 -125 1597 -115
rect 1492 -139 1496 -135
rect 1523 -139 1527 -135
rect 1554 -139 1558 -135
rect 1585 -139 1589 -135
rect 1486 -141 1589 -139
rect 1486 -145 1538 -141
rect 1542 -145 1589 -141
rect 1486 -151 1589 -149
rect 1486 -155 1540 -151
rect 1544 -155 1589 -151
rect 1231 -158 1235 -155
rect 1223 -163 1235 -158
rect 1282 -159 1286 -155
rect 1239 -163 1286 -159
rect 1492 -159 1496 -155
rect 1523 -159 1527 -155
rect 1554 -159 1558 -155
rect 1585 -159 1589 -155
rect 1225 -169 1249 -167
rect 1225 -173 1235 -169
rect 1239 -173 1249 -169
rect 1254 -173 1303 -167
rect 1231 -177 1235 -173
rect 1255 -177 1259 -173
rect 1299 -177 1303 -173
rect 1440 -191 1492 -186
rect 1515 -187 1519 -169
rect 1531 -180 1535 -169
rect 1562 -171 1566 -169
rect 1562 -175 1581 -171
rect 1531 -184 1555 -180
rect 1577 -184 1581 -175
rect 1593 -184 1597 -169
rect 1500 -191 1539 -187
rect 1239 -204 1243 -197
rect 1211 -208 1232 -204
rect 1239 -208 1256 -204
rect 1211 -234 1215 -208
rect 1239 -212 1243 -208
rect 1231 -226 1235 -222
rect 1223 -231 1235 -226
rect 1238 -230 1268 -226
rect 1238 -234 1242 -230
rect 1211 -238 1242 -234
rect 1245 -237 1270 -233
rect 1245 -242 1249 -237
rect 1277 -240 1281 -197
rect 1440 -240 1444 -191
rect 1500 -199 1504 -191
rect 1546 -199 1550 -184
rect 1577 -189 1585 -184
rect 1593 -189 1608 -184
rect 1577 -199 1581 -189
rect 1593 -199 1597 -189
rect 1492 -213 1496 -209
rect 1523 -213 1527 -209
rect 1554 -213 1558 -209
rect 1585 -213 1589 -209
rect 1486 -215 1589 -213
rect 1486 -219 1538 -215
rect 1542 -219 1589 -215
rect 1486 -225 1589 -223
rect 1486 -229 1540 -225
rect 1544 -229 1589 -225
rect 1218 -246 1249 -242
rect 1255 -244 1444 -240
rect 1492 -233 1496 -229
rect 1523 -233 1527 -229
rect 1554 -233 1558 -229
rect 1585 -233 1589 -229
rect 1218 -287 1222 -246
rect 1225 -252 1244 -250
rect 1225 -256 1235 -252
rect 1239 -256 1244 -252
rect 1231 -260 1235 -256
rect 1239 -287 1243 -280
rect 1069 -291 1232 -287
rect 1239 -292 1244 -287
rect 1239 -295 1243 -292
rect 1255 -295 1259 -244
rect 1263 -292 1297 -288
rect 1263 -295 1267 -292
rect 1293 -295 1297 -292
rect 1310 -295 1314 -244
rect 1439 -265 1492 -260
rect 1515 -261 1519 -243
rect 1531 -254 1535 -243
rect 1562 -245 1566 -243
rect 1562 -249 1581 -245
rect 1531 -258 1555 -254
rect 1577 -258 1581 -249
rect 1593 -258 1597 -243
rect 1500 -265 1539 -261
rect 1231 -308 1235 -305
rect 1223 -313 1235 -308
rect 1282 -309 1286 -305
rect 1239 -313 1286 -309
rect 1225 -319 1249 -317
rect 1225 -323 1235 -319
rect 1239 -323 1249 -319
rect 1254 -323 1303 -317
rect 1231 -327 1235 -323
rect 1255 -327 1259 -323
rect 1299 -327 1303 -323
rect 1239 -354 1243 -347
rect 1211 -358 1232 -354
rect 1239 -358 1256 -354
rect 1211 -384 1215 -358
rect 1239 -362 1243 -358
rect 1231 -376 1235 -372
rect 1223 -381 1235 -376
rect 1238 -380 1268 -376
rect 1238 -384 1242 -380
rect 1211 -388 1242 -384
rect 1245 -387 1270 -383
rect 1245 -392 1249 -387
rect 1277 -390 1281 -347
rect 1218 -396 1249 -392
rect 1255 -391 1314 -390
rect 1439 -391 1443 -265
rect 1500 -273 1504 -265
rect 1546 -273 1550 -258
rect 1577 -263 1585 -258
rect 1593 -263 1608 -258
rect 1577 -273 1581 -263
rect 1593 -273 1597 -263
rect 1492 -287 1496 -283
rect 1523 -287 1527 -283
rect 1554 -287 1558 -283
rect 1585 -287 1589 -283
rect 1486 -289 1589 -287
rect 1486 -293 1538 -289
rect 1542 -293 1589 -289
rect 1474 -303 1479 -301
rect 1486 -299 1589 -297
rect 1486 -303 1540 -299
rect 1544 -303 1589 -299
rect 1473 -306 1479 -303
rect 1473 -325 1478 -306
rect 1492 -307 1496 -303
rect 1523 -307 1527 -303
rect 1554 -307 1558 -303
rect 1585 -307 1589 -303
rect 1255 -394 1443 -391
rect 1218 -437 1222 -396
rect 1225 -402 1244 -400
rect 1225 -406 1235 -402
rect 1239 -406 1244 -402
rect 1231 -410 1235 -406
rect 1239 -437 1243 -430
rect 1019 -441 1232 -437
rect 1239 -442 1244 -437
rect 1239 -445 1243 -442
rect 1255 -445 1259 -394
rect 1310 -395 1443 -394
rect 1263 -442 1297 -438
rect 1263 -445 1267 -442
rect 1293 -445 1297 -442
rect 1310 -445 1314 -395
rect 1231 -458 1235 -455
rect 1223 -463 1235 -458
rect 1282 -459 1286 -455
rect 1239 -463 1286 -459
rect 796 -488 816 -482
rect 822 -484 1044 -482
rect 822 -488 844 -484
rect 848 -488 906 -484
rect 910 -488 968 -484
rect 972 -488 1030 -484
rect 1034 -488 1044 -484
rect 802 -492 806 -488
rect 840 -492 844 -488
rect 864 -492 868 -488
rect 902 -492 906 -488
rect 926 -492 930 -488
rect 964 -492 968 -488
rect 988 -492 992 -488
rect 1026 -492 1030 -488
rect 824 -519 828 -512
rect 848 -519 852 -512
rect 886 -519 890 -512
rect 910 -519 914 -512
rect 948 -519 952 -512
rect 972 -519 976 -512
rect 1010 -519 1014 -512
rect 1034 -519 1038 -512
rect 1454 -519 1458 -340
rect 748 -523 803 -519
rect 824 -523 841 -519
rect 848 -523 865 -519
rect 886 -523 903 -519
rect 910 -523 927 -519
rect 948 -523 965 -519
rect 972 -523 989 -519
rect 1010 -523 1027 -519
rect 1034 -523 1458 -519
rect 717 -530 817 -526
rect 246 -538 277 -534
rect 283 -536 479 -532
rect 246 -579 250 -538
rect 253 -544 272 -542
rect 253 -548 263 -544
rect 267 -548 272 -544
rect 259 -552 263 -548
rect 267 -579 271 -572
rect 242 -583 260 -579
rect 239 -646 243 -583
rect 267 -584 272 -579
rect 267 -587 271 -584
rect 283 -587 287 -536
rect 291 -584 325 -580
rect 291 -587 295 -584
rect 321 -587 325 -584
rect 338 -587 342 -536
rect 475 -537 479 -536
rect 505 -537 509 -530
rect 540 -537 544 -530
rect 567 -537 571 -530
rect 602 -537 606 -530
rect 824 -533 828 -523
rect 802 -537 828 -533
rect 475 -541 495 -537
rect 505 -541 533 -537
rect 540 -541 557 -537
rect 567 -541 595 -537
rect 602 -541 721 -537
rect 488 -548 509 -544
rect 516 -552 520 -541
rect 540 -552 544 -541
rect 554 -548 571 -544
rect 578 -552 582 -541
rect 602 -552 606 -541
rect 717 -562 721 -541
rect 802 -540 806 -537
rect 824 -540 828 -537
rect 848 -540 852 -523
rect 861 -530 879 -526
rect 886 -533 890 -523
rect 864 -537 890 -533
rect 864 -540 868 -537
rect 886 -540 890 -537
rect 910 -540 914 -523
rect 923 -530 941 -526
rect 948 -533 952 -523
rect 926 -537 952 -533
rect 926 -540 930 -537
rect 948 -540 952 -537
rect 972 -540 976 -523
rect 985 -530 1003 -526
rect 1010 -533 1014 -523
rect 988 -537 1014 -533
rect 988 -540 992 -537
rect 1010 -540 1014 -537
rect 1034 -540 1038 -523
rect 813 -554 817 -550
rect 840 -554 844 -550
rect 875 -554 879 -550
rect 902 -554 906 -550
rect 937 -554 941 -550
rect 964 -554 968 -550
rect 999 -554 1003 -550
rect 1026 -554 1030 -550
rect 799 -558 844 -554
rect 848 -558 906 -554
rect 910 -558 968 -554
rect 972 -558 1030 -554
rect 1034 -558 1039 -554
rect 494 -566 498 -562
rect 494 -570 504 -566
rect 532 -566 536 -562
rect 556 -566 560 -562
rect 594 -566 598 -562
rect 509 -570 536 -566
rect 540 -570 598 -566
rect 602 -570 612 -566
rect 717 -567 856 -562
rect 974 -567 980 -562
rect 544 -579 549 -574
rect 259 -600 263 -597
rect 251 -605 263 -600
rect 310 -601 314 -597
rect 267 -605 314 -601
rect 494 -602 545 -600
rect 494 -606 536 -602
rect 540 -606 545 -602
rect 249 -611 300 -609
rect 249 -615 291 -611
rect 295 -615 300 -611
rect 494 -610 498 -606
rect 516 -610 520 -606
rect 249 -619 253 -615
rect 271 -619 275 -615
rect 287 -619 291 -615
rect 532 -610 536 -606
rect 505 -637 509 -630
rect 540 -637 544 -630
rect 918 -637 923 -567
rect 260 -646 264 -639
rect 295 -646 299 -639
rect 488 -641 495 -637
rect 505 -641 533 -637
rect 540 -641 923 -637
rect 239 -650 250 -646
rect 260 -650 288 -646
rect 295 -650 351 -646
rect 488 -648 509 -644
rect 230 -657 264 -653
rect 271 -661 275 -650
rect 295 -661 299 -650
rect 516 -652 520 -641
rect 540 -652 544 -641
rect 494 -666 498 -662
rect 494 -670 504 -666
rect 532 -666 536 -662
rect 509 -670 536 -666
rect 540 -670 550 -666
rect 249 -674 253 -671
rect 251 -675 253 -674
rect 287 -675 291 -671
rect 251 -679 291 -675
rect 1473 -748 1478 -331
rect 1486 -335 1492 -334
rect 1489 -339 1492 -335
rect 1515 -335 1519 -317
rect 1531 -328 1535 -317
rect 1562 -319 1566 -317
rect 1562 -323 1581 -319
rect 1531 -332 1555 -328
rect 1577 -332 1581 -323
rect 1593 -332 1597 -317
rect 1500 -339 1539 -335
rect 1500 -347 1504 -339
rect 1546 -347 1550 -332
rect 1577 -337 1585 -332
rect 1593 -337 1608 -332
rect 1577 -347 1581 -337
rect 1593 -347 1597 -337
rect 1492 -361 1496 -357
rect 1523 -361 1527 -357
rect 1554 -361 1558 -357
rect 1585 -361 1589 -357
rect 1486 -363 1589 -361
rect 1486 -367 1538 -363
rect 1542 -367 1589 -363
rect -23 -753 1478 -748
<< m2contact >>
rect 607 251 612 257
rect 277 207 282 213
rect 326 207 331 213
rect 463 208 468 213
rect 246 149 251 154
rect 296 150 301 155
rect 3 36 8 41
rect 220 89 225 94
rect 3 -38 8 -33
rect 237 89 242 94
rect 272 124 277 130
rect 272 88 277 93
rect 487 208 492 213
rect 548 208 553 213
rect 504 186 509 191
rect 629 181 634 186
rect 548 172 553 177
rect 607 162 612 168
rect 246 67 251 72
rect 300 57 305 63
rect 246 -7 251 -2
rect 277 -17 282 -11
rect 326 -17 331 -11
rect 246 -75 251 -70
rect 296 -74 301 -69
rect 3 -112 8 -107
rect 220 -135 225 -130
rect 3 -186 8 -181
rect 486 118 491 123
rect 549 119 554 124
rect 504 98 509 103
rect 549 89 554 94
rect 641 116 647 122
rect 544 79 550 85
rect 691 73 696 78
rect 750 46 755 51
rect 691 37 696 42
rect 504 15 509 20
rect 616 -12 622 -6
rect 237 -135 242 -130
rect 272 -100 277 -94
rect 272 -136 277 -131
rect 246 -157 251 -152
rect 300 -167 305 -161
rect 246 -231 251 -226
rect 277 -241 282 -235
rect 326 -241 331 -235
rect 3 -260 8 -255
rect 246 -299 251 -294
rect 296 -298 301 -293
rect 3 -334 8 -329
rect 220 -359 225 -354
rect 3 -408 8 -403
rect 3 -482 8 -477
rect 237 -359 242 -354
rect 272 -324 277 -318
rect 272 -360 277 -355
rect 485 -56 490 -51
rect 548 -55 553 -50
rect 611 -55 616 -50
rect 504 -76 509 -71
rect 548 -85 553 -80
rect 611 -85 616 -80
rect 607 -109 612 -103
rect 719 -96 725 -90
rect 548 -152 553 -147
rect 778 -139 783 -134
rect 840 -139 845 -134
rect 504 -173 509 -168
rect 899 -166 904 -161
rect 778 -175 783 -170
rect 840 -175 845 -170
rect 548 -182 553 -177
rect 545 -194 550 -188
rect 504 -258 509 -253
rect 681 -306 687 -300
rect 486 -350 491 -344
rect 549 -349 554 -344
rect 610 -349 615 -344
rect 672 -349 677 -344
rect 504 -370 509 -365
rect 246 -381 251 -376
rect 549 -379 554 -374
rect 610 -379 615 -374
rect 672 -379 677 -374
rect 300 -391 305 -385
rect 669 -406 674 -400
rect 246 -455 251 -450
rect 549 -449 554 -444
rect 610 -449 615 -444
rect 277 -465 282 -459
rect 326 -465 331 -459
rect 504 -470 509 -465
rect 549 -479 554 -474
rect 610 -479 615 -474
rect 246 -523 251 -518
rect 296 -522 301 -517
rect 220 -583 225 -578
rect 607 -506 612 -500
rect 1249 127 1254 133
rect 1218 69 1223 74
rect 1268 70 1273 75
rect 1244 44 1249 50
rect 1244 8 1249 13
rect 1218 -13 1223 -8
rect 1249 -23 1254 -17
rect 1218 -81 1223 -76
rect 1268 -80 1273 -75
rect 1244 -106 1249 -100
rect 1244 -142 1249 -137
rect 1218 -163 1223 -158
rect 1249 -173 1254 -167
rect 1218 -231 1223 -226
rect 1268 -230 1273 -225
rect 1244 -256 1249 -250
rect 1244 -292 1249 -287
rect 1218 -313 1223 -308
rect 1249 -323 1254 -317
rect 1218 -381 1223 -376
rect 1268 -380 1273 -375
rect 1474 -301 1479 -296
rect 1473 -331 1479 -325
rect 1244 -406 1249 -400
rect 1244 -442 1249 -437
rect 1454 -340 1460 -334
rect 1218 -463 1223 -458
rect 816 -488 822 -482
rect 237 -583 242 -578
rect 272 -548 277 -542
rect 272 -584 277 -579
rect 549 -549 554 -544
rect 856 -531 861 -526
rect 918 -531 923 -526
rect 980 -531 985 -526
rect 1039 -558 1044 -553
rect 504 -570 509 -565
rect 856 -567 861 -562
rect 918 -567 923 -562
rect 980 -567 985 -562
rect 549 -579 554 -574
rect 246 -605 251 -600
rect 545 -606 550 -600
rect 300 -615 305 -609
rect 504 -670 509 -665
rect 246 -679 251 -674
rect 1483 -341 1489 -335
<< pm12contact >>
rect 21 36 26 41
rect 37 36 42 41
rect 83 36 88 41
rect 21 -38 26 -33
rect 37 -38 42 -33
rect 83 -38 88 -33
rect 319 150 324 155
rect 305 101 310 106
rect 21 -112 26 -107
rect 37 -112 42 -107
rect 83 -112 88 -107
rect 21 -186 26 -181
rect 37 -186 42 -181
rect 83 -186 88 -181
rect 319 -74 324 -69
rect 305 -123 310 -118
rect 21 -260 26 -255
rect 37 -260 42 -255
rect 83 -260 88 -255
rect 21 -334 26 -329
rect 37 -334 42 -329
rect 83 -334 88 -329
rect 21 -408 26 -403
rect 37 -408 42 -403
rect 83 -408 88 -403
rect 21 -482 26 -477
rect 37 -482 42 -477
rect 83 -482 88 -477
rect 319 -298 324 -293
rect 305 -347 310 -342
rect 319 -522 324 -517
rect 1291 70 1296 75
rect 1277 21 1282 26
rect 1507 -35 1512 -30
rect 1523 -35 1528 -30
rect 1569 -35 1574 -30
rect 1291 -80 1296 -75
rect 1277 -129 1282 -124
rect 1507 -109 1512 -104
rect 1523 -109 1528 -104
rect 1569 -109 1574 -104
rect 1507 -183 1512 -178
rect 1523 -183 1528 -178
rect 1569 -183 1574 -178
rect 1291 -230 1296 -225
rect 1277 -279 1282 -274
rect 1507 -257 1512 -252
rect 1523 -257 1528 -252
rect 1569 -257 1574 -252
rect 1291 -380 1296 -375
rect 1507 -331 1512 -326
rect 1277 -429 1282 -424
rect 305 -571 310 -566
rect 1523 -331 1528 -326
rect 1569 -331 1574 -326
<< ndm12contact >>
rect 299 75 304 85
rect 329 75 334 85
rect 299 -149 304 -139
rect 329 -149 334 -139
rect 299 -373 304 -363
rect 329 -373 334 -363
rect 1271 -5 1276 5
rect 1301 -5 1306 5
rect 1271 -155 1276 -145
rect 1301 -155 1306 -145
rect 1271 -305 1276 -295
rect 1301 -305 1306 -295
rect 1271 -455 1276 -445
rect 1301 -455 1306 -445
rect 299 -597 304 -587
rect 329 -597 334 -587
<< metal2 >>
rect 612 251 622 257
rect 331 207 347 213
rect 468 208 487 213
rect 225 89 237 94
rect 246 72 251 149
rect 277 124 282 207
rect 301 150 319 155
rect 277 101 305 106
rect 277 88 282 101
rect 299 88 334 92
rect 299 85 304 88
rect 329 85 334 88
rect 8 36 21 41
rect 26 36 37 41
rect 42 36 83 41
rect 246 -2 251 67
rect 341 63 347 207
rect 305 57 347 63
rect 8 -38 21 -33
rect 26 -38 37 -33
rect 42 -38 83 -33
rect 246 -70 251 -7
rect 341 -11 347 57
rect 8 -112 21 -107
rect 26 -112 37 -107
rect 42 -112 83 -107
rect 225 -135 237 -130
rect 246 -152 251 -75
rect 331 -17 347 -11
rect 277 -100 282 -17
rect 301 -74 319 -69
rect 277 -123 305 -118
rect 277 -136 282 -123
rect 299 -136 334 -132
rect 299 -139 304 -136
rect 329 -139 334 -136
rect 8 -186 21 -181
rect 26 -186 37 -181
rect 42 -186 83 -181
rect 246 -226 251 -157
rect 341 -161 347 -17
rect 305 -167 347 -161
rect 8 -260 21 -255
rect 26 -260 37 -255
rect 42 -260 83 -255
rect 246 -294 251 -231
rect 341 -235 347 -167
rect 8 -334 21 -329
rect 26 -334 37 -329
rect 42 -334 83 -329
rect 225 -359 237 -354
rect 246 -376 251 -299
rect 331 -241 347 -235
rect 277 -324 282 -241
rect 301 -298 319 -293
rect 277 -347 305 -342
rect 277 -360 282 -347
rect 299 -360 334 -356
rect 299 -363 304 -360
rect 329 -363 334 -360
rect 8 -408 21 -403
rect 26 -408 37 -403
rect 42 -408 83 -403
rect 246 -450 251 -381
rect 341 -385 347 -241
rect 473 123 478 208
rect 473 118 486 123
rect 473 -51 478 118
rect 504 103 509 186
rect 548 177 553 208
rect 616 168 622 251
rect 634 181 781 186
rect 612 162 647 168
rect 504 20 509 98
rect 549 94 554 119
rect 616 85 622 162
rect 641 122 647 162
rect 550 79 622 85
rect 473 -56 485 -51
rect 473 -345 478 -56
rect 504 -71 509 15
rect 616 11 622 79
rect 691 42 696 73
rect 776 51 781 181
rect 755 46 942 51
rect 616 5 725 11
rect 616 -6 622 5
rect 504 -168 509 -76
rect 548 -80 553 -55
rect 611 -80 616 -55
rect 719 -83 725 5
rect 681 -89 725 -83
rect 681 -103 687 -89
rect 719 -90 725 -89
rect 612 -109 687 -103
rect 504 -253 509 -173
rect 548 -177 553 -152
rect 681 -188 687 -109
rect 778 -170 783 -139
rect 840 -170 845 -139
rect 937 -159 942 46
rect 1218 -8 1223 69
rect 1249 44 1254 127
rect 1273 70 1291 75
rect 1249 21 1277 26
rect 1249 8 1254 21
rect 1271 8 1306 12
rect 1271 5 1276 8
rect 1301 5 1306 8
rect 1218 -158 1223 -81
rect 1249 -106 1254 -23
rect 1474 -35 1507 -30
rect 1512 -35 1523 -30
rect 1528 -35 1569 -30
rect 1273 -80 1291 -75
rect 1474 -104 1479 -35
rect 1474 -109 1507 -104
rect 1512 -109 1523 -104
rect 1528 -109 1569 -104
rect 1249 -129 1277 -124
rect 1249 -142 1254 -129
rect 1271 -142 1306 -138
rect 1271 -145 1276 -142
rect 1301 -145 1306 -142
rect 937 -161 1103 -159
rect 904 -164 1103 -161
rect 904 -166 942 -164
rect 550 -194 687 -188
rect 473 -350 486 -345
rect 305 -391 347 -385
rect 8 -482 21 -477
rect 26 -482 37 -477
rect 42 -482 83 -477
rect 246 -518 251 -455
rect 341 -459 347 -391
rect 225 -583 237 -578
rect 246 -600 251 -523
rect 331 -465 347 -459
rect 277 -548 282 -465
rect 301 -522 319 -517
rect 277 -571 305 -566
rect 277 -584 282 -571
rect 299 -584 334 -580
rect 299 -587 304 -584
rect 329 -587 334 -584
rect 246 -674 251 -605
rect 341 -609 347 -465
rect 305 -615 347 -609
rect 504 -365 509 -258
rect 681 -287 687 -194
rect 681 -293 822 -287
rect 681 -300 687 -293
rect 504 -465 509 -370
rect 549 -374 554 -349
rect 610 -374 615 -349
rect 672 -374 677 -349
rect 816 -400 822 -293
rect 674 -406 822 -400
rect 504 -565 509 -470
rect 549 -474 554 -449
rect 610 -474 615 -449
rect 697 -500 703 -406
rect 816 -482 822 -406
rect 612 -506 703 -500
rect 504 -665 509 -570
rect 549 -574 554 -549
rect 626 -600 632 -506
rect 856 -562 861 -531
rect 918 -562 923 -531
rect 980 -562 985 -531
rect 1098 -553 1103 -164
rect 1218 -308 1223 -231
rect 1249 -256 1254 -173
rect 1474 -178 1479 -109
rect 1474 -183 1507 -178
rect 1512 -183 1523 -178
rect 1528 -183 1569 -178
rect 1273 -230 1291 -225
rect 1474 -252 1479 -183
rect 1474 -257 1507 -252
rect 1512 -257 1523 -252
rect 1528 -257 1569 -252
rect 1249 -279 1277 -274
rect 1249 -292 1254 -279
rect 1271 -292 1306 -288
rect 1271 -295 1276 -292
rect 1301 -295 1306 -292
rect 1474 -296 1479 -257
rect 1218 -458 1223 -381
rect 1249 -406 1254 -323
rect 1479 -331 1507 -326
rect 1512 -331 1523 -326
rect 1528 -331 1569 -326
rect 1460 -340 1483 -335
rect 1454 -341 1483 -340
rect 1273 -380 1291 -375
rect 1249 -429 1277 -424
rect 1249 -442 1254 -429
rect 1271 -442 1306 -438
rect 1271 -445 1276 -442
rect 1301 -445 1306 -442
rect 1044 -558 1103 -553
rect 550 -606 632 -600
<< labels >>
rlabel metal1 2 3 2 3 2 gnd
rlabel metal1 2 67 2 67 4 vdd
rlabel metal1 2 -71 2 -71 2 gnd
rlabel metal1 2 -7 2 -7 4 vdd
rlabel metal1 2 -145 2 -145 2 gnd
rlabel metal1 2 -81 2 -81 4 vdd
rlabel metal1 2 -219 2 -219 2 gnd
rlabel metal1 2 -155 2 -155 4 vdd
rlabel metal1 2 -293 2 -293 2 gnd
rlabel metal1 2 -229 2 -229 4 vdd
rlabel metal1 2 -367 2 -367 2 gnd
rlabel metal1 2 -303 2 -303 4 vdd
rlabel metal1 2 -441 2 -441 2 gnd
rlabel metal1 2 -377 2 -377 4 vdd
rlabel metal1 2 -515 2 -515 2 gnd
rlabel metal1 2 -451 2 -451 4 vdd
rlabel metal1 255 210 255 210 5 vdd
rlabel metal1 350 138 350 138 7 P0
rlabel metal1 350 24 350 24 7 G0
rlabel metal1 350 -86 350 -86 7 P1
rlabel metal1 350 -200 350 -200 7 G1
rlabel metal1 350 -310 350 -310 7 P2
rlabel metal1 350 -424 350 -424 7 G2
rlabel metal1 350 -534 350 -534 7 P3
rlabel metal1 349 -648 349 -648 7 G3
rlabel metal1 274 -677 274 -677 1 gnd
rlabel metal1 610 218 610 218 1 C1
rlabel metal1 754 83 754 83 7 C2
rlabel metal1 903 -129 903 -129 1 C3
rlabel metal1 1042 -521 1042 -521 7 Cout
rlabel metal1 523 -668 523 -668 1 gnd
rlabel metal1 549 254 549 254 5 vdd
rlabel metal1 475 218 475 218 3 Cin
rlabel metal1 459 210 459 210 3 P0
rlabel metal1 491 174 491 174 1 G0
rlabel metal1 488 91 488 91 1 P1
rlabel metal1 490 39 490 39 1 G0
rlabel metal1 662 39 662 39 1 G1
rlabel metal1 604 -83 604 -83 1 P2
rlabel metal1 540 -83 540 -83 1 P1
rlabel metal1 491 -149 491 -149 1 P2
rlabel metal1 542 -180 542 -180 1 G0
rlabel metal1 490 -227 490 -227 1 P2
rlabel metal1 490 -234 490 -234 1 G1
rlabel metal1 835 -173 835 -173 1 G2
rlabel metal1 546 -377 546 -377 1 P1
rlabel metal1 490 -439 490 -439 1 P1
rlabel metal1 606 -376 606 -376 1 P2
rlabel metal1 490 -446 490 -446 1 P2
rlabel metal1 667 -377 667 -377 1 P3
rlabel metal1 545 -477 545 -477 1 P3
rlabel metal1 605 -477 605 -477 1 G0
rlabel metal1 490 -539 490 -539 1 P3
rlabel metal1 490 -546 490 -546 1 P2
rlabel metal1 546 -577 546 -577 1 G1
rlabel metal1 489 -639 489 -639 1 P3
rlabel metal1 489 -646 489 -646 1 G2
rlabel metal1 976 -565 976 -565 1 G3
rlabel metal1 1228 130 1228 130 4 vdd
rlabel metal1 1227 -11 1227 -11 2 gnd
rlabel metal1 1312 58 1312 58 7 S0
rlabel metal1 1226 94 1226 94 1 P0
rlabel metal1 1226 11 1226 11 1 Cin
rlabel metal1 1228 -20 1228 -20 4 vdd
rlabel metal1 1227 -161 1227 -161 2 gnd
rlabel metal1 1228 -170 1228 -170 4 vdd
rlabel metal1 1227 -311 1227 -311 2 gnd
rlabel metal1 1228 -320 1228 -320 4 vdd
rlabel metal1 1227 -461 1227 -461 2 gnd
rlabel metal1 1226 -56 1226 -56 1 P1
rlabel metal1 1226 -139 1226 -139 1 C1
rlabel metal1 1226 -206 1226 -206 1 P2
rlabel metal1 1226 -289 1226 -289 1 C2
rlabel metal1 1226 -356 1226 -356 1 P3
rlabel metal1 1226 -439 1226 -439 1 C3
rlabel metal1 1312 -392 1312 -392 7 S3
rlabel metal1 1312 -242 1312 -242 7 S2
rlabel metal1 1312 -92 1312 -92 7 S1
rlabel metal1 1488 -4 1488 -4 4 vdd
rlabel metal1 1488 -290 1488 -290 2 gnd
rlabel metal1 1 30 1 30 3 A0
rlabel metal1 1 -44 1 -44 3 B0
rlabel metal1 1 -118 1 -118 3 A1
rlabel metal1 1 -192 1 -192 3 B1
rlabel metal1 1 -266 1 -266 3 A2
rlabel metal1 1 -340 1 -340 3 B2
rlabel metal1 1 -414 1 -414 3 A3
rlabel metal1 1 -488 1 -488 3 B3
rlabel metal1 -20 -533 -20 -533 3 clk
rlabel metal1 1606 -39 1606 -39 7 S0
rlabel metal1 1606 -113 1606 -113 7 S1
rlabel metal1 1606 -187 1606 -187 7 S2
rlabel metal1 1606 -261 1606 -261 7 S3
rlabel metal1 1488 -364 1488 -364 2 gnd
rlabel metal1 1606 -335 1606 -335 7 Cout
<< end >>
