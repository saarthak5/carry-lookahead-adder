* Propagate & Generate

.include TSMC_180nm.txt
.param SUPPLY=1.8
.param LAMBDA=0.09u
.param Wn={10*LAMBDA}
.param Wp={2*Wn}
.global gnd vdd

* Source		Nodes			Value
*****************************************
Vdd				vdd	gnd			'SUPPLY'
Va0				a0	gnd			'SUPPLY'
Va1				a1	gnd			'SUPPLY'
Va2				a2	gnd			'SUPPLY'
Va3				a3	gnd				0
Vb0				b0	gnd				0
Vb1				b1	gnd			'SUPPLY'
Vb2				b2	gnd				0
Vb3				b3	gnd			'SUPPLY'

* A = 0111, B = 1010

.subckt INV x xbar

Mp xbar x vdd vdd CMOSP
+ L={2*LAMBDA} W={Wp}
+ AS={5*Wp*LAMBDA} AD={5*Wp*LAMBDA}
+ PS={10*LAMBDA+2*Wp} PD={10*LAMBDA+2*Wp}

Mn xbar x gnd gnd CMOSN
+ L={2*LAMBDA} W={Wn}
+ AS={5*Wn*LAMBDA} AD={5*Wn*LAMBDA}
+ PS={10*LAMBDA+2*Wn} PD={10*LAMBDA+2*Wn}

.ends INV

.subckt XOR f x y

X1 x xbar INV
X2 y ybar INV

Mp1 n1 x vdd vdd CMOSP
+ L={2*LAMBDA} W={Wp}
+ AS={5*Wp*LAMBDA} AD={5*Wp*LAMBDA}
+ PS={10*LAMBDA+2*Wp} PD={10*LAMBDA+2*Wp}

Mp2 n2 xbar vdd vdd CMOSP
+ L={2*LAMBDA} W={Wp}
+ AS={5*Wp*LAMBDA} AD={5*Wp*LAMBDA}
+ PS={10*LAMBDA+2*Wp} PD={10*LAMBDA+2*Wp}

Mp3 f ybar n1 vdd CMOSP
+ L={2*LAMBDA} W={Wp}
+ AS={5*Wp*LAMBDA} AD={5*Wp*LAMBDA}
+ PS={10*LAMBDA+2*Wp} PD={10*LAMBDA+2*Wp}

Mp4 f y n2 vdd CMOSP
+ L={2*LAMBDA} W={Wp}
+ AS={5*Wp*LAMBDA} AD={5*Wp*LAMBDA}
+ PS={10*LAMBDA+2*Wp} PD={10*LAMBDA+2*Wp}

Mn1 f xbar n3 gnd CMOSN
+ L={2*LAMBDA} W={Wn}
+ AS={5*Wn*LAMBDA} AD={5*Wn*LAMBDA}
+ PS={10*LAMBDA+2*Wn} PD={10*LAMBDA+2*Wn}

Mn2 f x n4 gnd CMOSN
+ L={2*LAMBDA} W={Wn}
+ AS={5*Wn*LAMBDA} AD={5*Wn*LAMBDA}
+ PS={10*LAMBDA+2*Wn} PD={10*LAMBDA+2*Wn}

Mn3 n3 ybar gnd gnd CMOSN
+ L={2*LAMBDA} W={Wn}
+ AS={5*Wn*LAMBDA} AD={5*Wn*LAMBDA}
+ PS={10*LAMBDA+2*Wn} PD={10*LAMBDA+2*Wn}

Mn4 n4 y gnd gnd CMOSN
+ L={2*LAMBDA} W={Wn}
+ AS={5*Wn*LAMBDA} AD={5*Wn*LAMBDA}
+ PS={10*LAMBDA+2*Wn} PD={10*LAMBDA+2*Wn}

.ends XOR

.subckt AND f x y

.param Wp={2*Wn}
Mp1 fbar x vdd vdd CMOSP
+ L={2*LAMBDA} W={Wp}
+ AS={5*Wp*LAMBDA} AD={5*Wp*LAMBDA}
+ PS={10*LAMBDA+2*Wp} PD={10*LAMBDA+2*Wp}

Mp2 fbar y vdd vdd CMOSP
+ L={2*LAMBDA} W={Wp}
+ AS={5*Wp*LAMBDA} AD={5*Wp*LAMBDA}
+ PS={10*LAMBDA+2*Wp} PD={10*LAMBDA+2*Wp}

Mn1 fbar x n1 gnd CMOSN
+ L={2*LAMBDA} W={Wn}
+ AS={5*Wn*LAMBDA} AD={5*Wn*LAMBDA}
+ PS={10*LAMBDA+2*Wn} PD={10*LAMBDA+2*Wn}

Mn2 n1 y gnd gnd CMOSN
+ L={2*LAMBDA} W={Wn}
+ AS={5*Wn*LAMBDA} AD={5*Wn*LAMBDA}
+ PS={10*LAMBDA+2*Wn} PD={10*LAMBDA+2*Wn}

X1 fbar f INV

.ends AND

.subckt PG p0 p1 p2 p3 g0 g1 g2 g3 a0 a1 a2 a3 b0 b1 b2 b3

Xp0 p0 a0 b0 XOR
Xp1 p1 a1 b1 XOR
Xp2 p2 a2 b2 XOR
Xp3 p3 a3 b3 XOR

Xg0 g0 a0 b0 AND
Xg1 g1 a1 b1 AND
Xg2 g2 a2 b2 AND
Xg3 g3 a3 b3 AND

.ends PG

X1 p0 p1 p2 p3 g0 g1 g2 g3 a0 a1 a2 a3 b0 b1 b2 b3 PG

.control
tran 10p 20p
run

set hcopypscolor=1
set color0=white
set color1=black

plot V(p0) V(p1)+2 V(p2)+4 V(p3)+6 V(g0)+8 V(g1)+10 V(g2)+12 V(g3)+14
hardcopy V(p0) V(p1)+2 V(p2)+4 V(p3)+6 V(g0)+8 V(g1)+10 V(g2)+12 V(g3)+14
.endc

.end
