magic
tech scmos
timestamp 1732088497
<< nwell >>
rect 0 34 124 71
rect 0 -55 124 -18
rect 143 -101 267 -64
rect 0 -138 62 -101
rect 0 -229 186 -192
rect 0 -326 124 -289
rect 230 -313 416 -276
rect 0 -411 62 -374
rect 0 -523 248 -486
rect 0 -623 186 -586
rect 0 -723 124 -686
rect 308 -705 556 -668
rect 0 -823 62 -786
<< ntransistor >>
rect 11 8 13 18
rect 25 8 27 18
rect 49 8 51 18
rect 73 2 75 12
rect 87 2 89 12
rect 111 2 113 12
rect 11 -81 13 -71
rect 25 -81 27 -71
rect 49 -81 51 -71
rect 73 -81 75 -71
rect 87 -81 89 -71
rect 111 -81 113 -71
rect 154 -133 156 -123
rect 168 -133 170 -123
rect 192 -133 194 -123
rect 216 -133 218 -123
rect 230 -133 232 -123
rect 254 -133 256 -123
rect 11 -164 13 -154
rect 25 -164 27 -154
rect 49 -164 51 -154
rect 11 -255 13 -245
rect 25 -255 27 -245
rect 49 -255 51 -245
rect 73 -255 75 -245
rect 87 -255 89 -245
rect 111 -255 113 -245
rect 135 -255 137 -245
rect 149 -255 151 -245
rect 173 -255 175 -245
rect 11 -352 13 -342
rect 25 -352 27 -342
rect 49 -352 51 -342
rect 73 -352 75 -342
rect 87 -352 89 -342
rect 111 -352 113 -342
rect 241 -345 243 -335
rect 255 -345 257 -335
rect 279 -345 281 -335
rect 303 -345 305 -335
rect 317 -345 319 -335
rect 341 -345 343 -335
rect 365 -345 367 -335
rect 379 -345 381 -335
rect 403 -345 405 -335
rect 11 -437 13 -427
rect 25 -437 27 -427
rect 49 -437 51 -427
rect 11 -549 13 -539
rect 25 -549 27 -539
rect 49 -549 51 -539
rect 73 -549 75 -539
rect 87 -549 89 -539
rect 111 -549 113 -539
rect 135 -549 137 -539
rect 149 -549 151 -539
rect 173 -549 175 -539
rect 197 -549 199 -539
rect 211 -549 213 -539
rect 235 -549 237 -539
rect 11 -649 13 -639
rect 25 -649 27 -639
rect 49 -649 51 -639
rect 73 -649 75 -639
rect 87 -649 89 -639
rect 111 -649 113 -639
rect 135 -649 137 -639
rect 149 -649 151 -639
rect 173 -649 175 -639
rect 319 -737 321 -727
rect 333 -737 335 -727
rect 357 -737 359 -727
rect 381 -737 383 -727
rect 395 -737 397 -727
rect 419 -737 421 -727
rect 443 -737 445 -727
rect 457 -737 459 -727
rect 481 -737 483 -727
rect 505 -737 507 -727
rect 519 -737 521 -727
rect 543 -737 545 -727
rect 11 -749 13 -739
rect 25 -749 27 -739
rect 49 -749 51 -739
rect 73 -749 75 -739
rect 87 -749 89 -739
rect 111 -749 113 -739
rect 11 -849 13 -839
rect 25 -849 27 -839
rect 49 -849 51 -839
<< ptransistor >>
rect 11 40 13 60
rect 25 40 27 60
rect 49 40 51 60
rect 73 40 75 60
rect 87 40 89 60
rect 111 40 113 60
rect 11 -49 13 -29
rect 25 -49 27 -29
rect 49 -49 51 -29
rect 73 -49 75 -29
rect 87 -49 89 -29
rect 111 -49 113 -29
rect 154 -95 156 -75
rect 168 -95 170 -75
rect 192 -95 194 -75
rect 216 -95 218 -75
rect 230 -95 232 -75
rect 254 -95 256 -75
rect 11 -132 13 -112
rect 25 -132 27 -112
rect 49 -132 51 -112
rect 11 -223 13 -203
rect 25 -223 27 -203
rect 49 -223 51 -203
rect 73 -223 75 -203
rect 87 -223 89 -203
rect 111 -223 113 -203
rect 135 -223 137 -203
rect 149 -223 151 -203
rect 173 -223 175 -203
rect 11 -320 13 -300
rect 25 -320 27 -300
rect 49 -320 51 -300
rect 73 -320 75 -300
rect 87 -320 89 -300
rect 111 -320 113 -300
rect 241 -307 243 -287
rect 255 -307 257 -287
rect 279 -307 281 -287
rect 303 -307 305 -287
rect 317 -307 319 -287
rect 341 -307 343 -287
rect 365 -307 367 -287
rect 379 -307 381 -287
rect 403 -307 405 -287
rect 11 -405 13 -385
rect 25 -405 27 -385
rect 49 -405 51 -385
rect 11 -517 13 -497
rect 25 -517 27 -497
rect 49 -517 51 -497
rect 73 -517 75 -497
rect 87 -517 89 -497
rect 111 -517 113 -497
rect 135 -517 137 -497
rect 149 -517 151 -497
rect 173 -517 175 -497
rect 197 -517 199 -497
rect 211 -517 213 -497
rect 235 -517 237 -497
rect 11 -617 13 -597
rect 25 -617 27 -597
rect 49 -617 51 -597
rect 73 -617 75 -597
rect 87 -617 89 -597
rect 111 -617 113 -597
rect 135 -617 137 -597
rect 149 -617 151 -597
rect 173 -617 175 -597
rect 11 -717 13 -697
rect 25 -717 27 -697
rect 49 -717 51 -697
rect 73 -717 75 -697
rect 87 -717 89 -697
rect 111 -717 113 -697
rect 319 -699 321 -679
rect 333 -699 335 -679
rect 357 -699 359 -679
rect 381 -699 383 -679
rect 395 -699 397 -679
rect 419 -699 421 -679
rect 443 -699 445 -679
rect 457 -699 459 -679
rect 481 -699 483 -679
rect 505 -699 507 -679
rect 519 -699 521 -679
rect 543 -699 545 -679
rect 11 -817 13 -797
rect 25 -817 27 -797
rect 49 -817 51 -797
<< ndiffusion >>
rect 10 8 11 18
rect 13 8 25 18
rect 27 8 28 18
rect 48 8 49 18
rect 51 8 52 18
rect 72 2 73 12
rect 75 2 79 12
rect 83 2 87 12
rect 89 2 90 12
rect 110 2 111 12
rect 113 2 114 12
rect 10 -81 11 -71
rect 13 -81 25 -71
rect 27 -81 28 -71
rect 48 -81 49 -71
rect 51 -81 52 -71
rect 72 -81 73 -71
rect 75 -81 87 -71
rect 89 -81 90 -71
rect 110 -81 111 -71
rect 113 -81 114 -71
rect 153 -133 154 -123
rect 156 -133 160 -123
rect 164 -133 168 -123
rect 170 -133 171 -123
rect 191 -133 192 -123
rect 194 -133 195 -123
rect 215 -133 216 -123
rect 218 -133 222 -123
rect 226 -133 230 -123
rect 232 -133 233 -123
rect 253 -133 254 -123
rect 256 -133 257 -123
rect 10 -164 11 -154
rect 13 -164 25 -154
rect 27 -164 28 -154
rect 48 -164 49 -154
rect 51 -164 52 -154
rect 10 -255 11 -245
rect 13 -255 25 -245
rect 27 -255 28 -245
rect 48 -255 49 -245
rect 51 -255 52 -245
rect 72 -255 73 -245
rect 75 -255 87 -245
rect 89 -255 90 -245
rect 110 -255 111 -245
rect 113 -255 114 -245
rect 134 -255 135 -245
rect 137 -255 149 -245
rect 151 -255 152 -245
rect 172 -255 173 -245
rect 175 -255 176 -245
rect 10 -352 11 -342
rect 13 -352 25 -342
rect 27 -352 28 -342
rect 48 -352 49 -342
rect 51 -352 52 -342
rect 72 -352 73 -342
rect 75 -352 87 -342
rect 89 -352 90 -342
rect 110 -352 111 -342
rect 113 -352 114 -342
rect 240 -345 241 -335
rect 243 -345 247 -335
rect 251 -345 255 -335
rect 257 -345 258 -335
rect 278 -345 279 -335
rect 281 -345 282 -335
rect 302 -345 303 -335
rect 305 -345 309 -335
rect 313 -345 317 -335
rect 319 -345 320 -335
rect 340 -345 341 -335
rect 343 -345 344 -335
rect 364 -345 365 -335
rect 367 -345 371 -335
rect 375 -345 379 -335
rect 381 -345 382 -335
rect 402 -345 403 -335
rect 405 -345 406 -335
rect 10 -437 11 -427
rect 13 -437 25 -427
rect 27 -437 28 -427
rect 48 -437 49 -427
rect 51 -437 52 -427
rect 10 -549 11 -539
rect 13 -549 25 -539
rect 27 -549 28 -539
rect 48 -549 49 -539
rect 51 -549 52 -539
rect 72 -549 73 -539
rect 75 -549 87 -539
rect 89 -549 90 -539
rect 110 -549 111 -539
rect 113 -549 114 -539
rect 134 -549 135 -539
rect 137 -549 149 -539
rect 151 -549 152 -539
rect 172 -549 173 -539
rect 175 -549 176 -539
rect 196 -549 197 -539
rect 199 -549 211 -539
rect 213 -549 214 -539
rect 234 -549 235 -539
rect 237 -549 238 -539
rect 10 -649 11 -639
rect 13 -649 25 -639
rect 27 -649 28 -639
rect 48 -649 49 -639
rect 51 -649 52 -639
rect 72 -649 73 -639
rect 75 -649 87 -639
rect 89 -649 90 -639
rect 110 -649 111 -639
rect 113 -649 114 -639
rect 134 -649 135 -639
rect 137 -649 149 -639
rect 151 -649 152 -639
rect 172 -649 173 -639
rect 175 -649 176 -639
rect 318 -737 319 -727
rect 321 -737 325 -727
rect 329 -737 333 -727
rect 335 -737 336 -727
rect 356 -737 357 -727
rect 359 -737 360 -727
rect 380 -737 381 -727
rect 383 -737 387 -727
rect 391 -737 395 -727
rect 397 -737 398 -727
rect 418 -737 419 -727
rect 421 -737 422 -727
rect 442 -737 443 -727
rect 445 -737 449 -727
rect 453 -737 457 -727
rect 459 -737 460 -727
rect 480 -737 481 -727
rect 483 -737 484 -727
rect 504 -737 505 -727
rect 507 -737 511 -727
rect 515 -737 519 -727
rect 521 -737 522 -727
rect 542 -737 543 -727
rect 545 -737 546 -727
rect 10 -749 11 -739
rect 13 -749 25 -739
rect 27 -749 28 -739
rect 48 -749 49 -739
rect 51 -749 52 -739
rect 72 -749 73 -739
rect 75 -749 87 -739
rect 89 -749 90 -739
rect 110 -749 111 -739
rect 113 -749 114 -739
rect 10 -849 11 -839
rect 13 -849 25 -839
rect 27 -849 28 -839
rect 48 -849 49 -839
rect 51 -849 52 -839
<< pdiffusion >>
rect 10 40 11 60
rect 13 40 17 60
rect 21 40 25 60
rect 27 40 28 60
rect 48 40 49 60
rect 51 40 52 60
rect 72 40 73 60
rect 75 40 87 60
rect 89 40 90 60
rect 110 40 111 60
rect 113 40 114 60
rect 10 -49 11 -29
rect 13 -49 17 -29
rect 21 -49 25 -29
rect 27 -49 28 -29
rect 48 -49 49 -29
rect 51 -49 52 -29
rect 72 -49 73 -29
rect 75 -49 79 -29
rect 83 -49 87 -29
rect 89 -49 90 -29
rect 110 -49 111 -29
rect 113 -49 114 -29
rect 153 -95 154 -75
rect 156 -95 168 -75
rect 170 -95 171 -75
rect 191 -95 192 -75
rect 194 -95 195 -75
rect 215 -95 216 -75
rect 218 -95 230 -75
rect 232 -95 233 -75
rect 253 -95 254 -75
rect 256 -95 257 -75
rect 10 -132 11 -112
rect 13 -132 17 -112
rect 21 -132 25 -112
rect 27 -132 28 -112
rect 48 -132 49 -112
rect 51 -132 52 -112
rect 10 -223 11 -203
rect 13 -223 17 -203
rect 21 -223 25 -203
rect 27 -223 28 -203
rect 48 -223 49 -203
rect 51 -223 52 -203
rect 72 -223 73 -203
rect 75 -223 79 -203
rect 83 -223 87 -203
rect 89 -223 90 -203
rect 110 -223 111 -203
rect 113 -223 114 -203
rect 134 -223 135 -203
rect 137 -223 141 -203
rect 145 -223 149 -203
rect 151 -223 152 -203
rect 172 -223 173 -203
rect 175 -223 176 -203
rect 10 -320 11 -300
rect 13 -320 17 -300
rect 21 -320 25 -300
rect 27 -320 28 -300
rect 48 -320 49 -300
rect 51 -320 52 -300
rect 72 -320 73 -300
rect 75 -320 79 -300
rect 83 -320 87 -300
rect 89 -320 90 -300
rect 110 -320 111 -300
rect 113 -320 114 -300
rect 240 -307 241 -287
rect 243 -307 255 -287
rect 257 -307 258 -287
rect 278 -307 279 -287
rect 281 -307 282 -287
rect 302 -307 303 -287
rect 305 -307 317 -287
rect 319 -307 320 -287
rect 340 -307 341 -287
rect 343 -307 344 -287
rect 364 -307 365 -287
rect 367 -307 379 -287
rect 381 -307 382 -287
rect 402 -307 403 -287
rect 405 -307 406 -287
rect 10 -405 11 -385
rect 13 -405 17 -385
rect 21 -405 25 -385
rect 27 -405 28 -385
rect 48 -405 49 -385
rect 51 -405 52 -385
rect 10 -517 11 -497
rect 13 -517 17 -497
rect 21 -517 25 -497
rect 27 -517 28 -497
rect 48 -517 49 -497
rect 51 -517 52 -497
rect 72 -517 73 -497
rect 75 -517 79 -497
rect 83 -517 87 -497
rect 89 -517 90 -497
rect 110 -517 111 -497
rect 113 -517 114 -497
rect 134 -517 135 -497
rect 137 -517 141 -497
rect 145 -517 149 -497
rect 151 -517 152 -497
rect 172 -517 173 -497
rect 175 -517 176 -497
rect 196 -517 197 -497
rect 199 -517 203 -497
rect 207 -517 211 -497
rect 213 -517 214 -497
rect 234 -517 235 -497
rect 237 -517 238 -497
rect 10 -617 11 -597
rect 13 -617 17 -597
rect 21 -617 25 -597
rect 27 -617 28 -597
rect 48 -617 49 -597
rect 51 -617 52 -597
rect 72 -617 73 -597
rect 75 -617 79 -597
rect 83 -617 87 -597
rect 89 -617 90 -597
rect 110 -617 111 -597
rect 113 -617 114 -597
rect 134 -617 135 -597
rect 137 -617 141 -597
rect 145 -617 149 -597
rect 151 -617 152 -597
rect 172 -617 173 -597
rect 175 -617 176 -597
rect 10 -717 11 -697
rect 13 -717 17 -697
rect 21 -717 25 -697
rect 27 -717 28 -697
rect 48 -717 49 -697
rect 51 -717 52 -697
rect 72 -717 73 -697
rect 75 -717 79 -697
rect 83 -717 87 -697
rect 89 -717 90 -697
rect 110 -717 111 -697
rect 113 -717 114 -697
rect 318 -699 319 -679
rect 321 -699 333 -679
rect 335 -699 336 -679
rect 356 -699 357 -679
rect 359 -699 360 -679
rect 380 -699 381 -679
rect 383 -699 395 -679
rect 397 -699 398 -679
rect 418 -699 419 -679
rect 421 -699 422 -679
rect 442 -699 443 -679
rect 445 -699 457 -679
rect 459 -699 460 -679
rect 480 -699 481 -679
rect 483 -699 484 -679
rect 504 -699 505 -679
rect 507 -699 519 -679
rect 521 -699 522 -679
rect 542 -699 543 -679
rect 545 -699 546 -679
rect 10 -817 11 -797
rect 13 -817 17 -797
rect 21 -817 25 -797
rect 27 -817 28 -797
rect 48 -817 49 -797
rect 51 -817 52 -797
<< ndcontact >>
rect 6 8 10 18
rect 28 8 32 18
rect 44 8 48 18
rect 52 8 56 18
rect 68 2 72 12
rect 79 2 83 12
rect 90 2 94 12
rect 106 2 110 12
rect 114 2 118 12
rect 6 -81 10 -71
rect 28 -81 32 -71
rect 44 -81 48 -71
rect 52 -81 56 -71
rect 68 -81 72 -71
rect 90 -81 94 -71
rect 106 -81 110 -71
rect 114 -81 118 -71
rect 149 -133 153 -123
rect 160 -133 164 -123
rect 171 -133 175 -123
rect 187 -133 191 -123
rect 195 -133 199 -123
rect 211 -133 215 -123
rect 222 -133 226 -123
rect 233 -133 237 -123
rect 249 -133 253 -123
rect 257 -133 261 -123
rect 6 -164 10 -154
rect 28 -164 32 -154
rect 44 -164 48 -154
rect 52 -164 56 -154
rect 6 -255 10 -245
rect 28 -255 32 -245
rect 44 -255 48 -245
rect 52 -255 56 -245
rect 68 -255 72 -245
rect 90 -255 94 -245
rect 106 -255 110 -245
rect 114 -255 118 -245
rect 130 -255 134 -245
rect 152 -255 156 -245
rect 168 -255 172 -245
rect 176 -255 180 -245
rect 6 -352 10 -342
rect 28 -352 32 -342
rect 44 -352 48 -342
rect 52 -352 56 -342
rect 68 -352 72 -342
rect 90 -352 94 -342
rect 106 -352 110 -342
rect 114 -352 118 -342
rect 236 -345 240 -335
rect 247 -345 251 -335
rect 258 -345 262 -335
rect 274 -345 278 -335
rect 282 -345 286 -335
rect 298 -345 302 -335
rect 309 -345 313 -335
rect 320 -345 324 -335
rect 336 -345 340 -335
rect 344 -345 348 -335
rect 360 -345 364 -335
rect 371 -345 375 -335
rect 382 -345 386 -335
rect 398 -345 402 -335
rect 406 -345 410 -335
rect 6 -437 10 -427
rect 28 -437 32 -427
rect 44 -437 48 -427
rect 52 -437 56 -427
rect 6 -549 10 -539
rect 28 -549 32 -539
rect 44 -549 48 -539
rect 52 -549 56 -539
rect 68 -549 72 -539
rect 90 -549 94 -539
rect 106 -549 110 -539
rect 114 -549 118 -539
rect 130 -549 134 -539
rect 152 -549 156 -539
rect 168 -549 172 -539
rect 176 -549 180 -539
rect 192 -549 196 -539
rect 214 -549 218 -539
rect 230 -549 234 -539
rect 238 -549 242 -539
rect 6 -649 10 -639
rect 28 -649 32 -639
rect 44 -649 48 -639
rect 52 -649 56 -639
rect 68 -649 72 -639
rect 90 -649 94 -639
rect 106 -649 110 -639
rect 114 -649 118 -639
rect 130 -649 134 -639
rect 152 -649 156 -639
rect 168 -649 172 -639
rect 176 -649 180 -639
rect 314 -737 318 -727
rect 325 -737 329 -727
rect 336 -737 340 -727
rect 352 -737 356 -727
rect 360 -737 364 -727
rect 376 -737 380 -727
rect 387 -737 391 -727
rect 398 -737 402 -727
rect 414 -737 418 -727
rect 422 -737 426 -727
rect 438 -737 442 -727
rect 449 -737 453 -727
rect 460 -737 464 -727
rect 476 -737 480 -727
rect 484 -737 488 -727
rect 500 -737 504 -727
rect 511 -737 515 -727
rect 522 -737 526 -727
rect 538 -737 542 -727
rect 546 -737 550 -727
rect 6 -749 10 -739
rect 28 -749 32 -739
rect 44 -749 48 -739
rect 52 -749 56 -739
rect 68 -749 72 -739
rect 90 -749 94 -739
rect 106 -749 110 -739
rect 114 -749 118 -739
rect 6 -849 10 -839
rect 28 -849 32 -839
rect 44 -849 48 -839
rect 52 -849 56 -839
<< pdcontact >>
rect 6 40 10 60
rect 17 40 21 60
rect 28 40 32 60
rect 44 40 48 60
rect 52 40 56 60
rect 68 40 72 60
rect 90 40 94 60
rect 106 40 110 60
rect 114 40 118 60
rect 6 -49 10 -29
rect 17 -49 21 -29
rect 28 -49 32 -29
rect 44 -49 48 -29
rect 52 -49 56 -29
rect 68 -49 72 -29
rect 79 -49 83 -29
rect 90 -49 94 -29
rect 106 -49 110 -29
rect 114 -49 118 -29
rect 149 -95 153 -75
rect 171 -95 175 -75
rect 187 -95 191 -75
rect 195 -95 199 -75
rect 211 -95 215 -75
rect 233 -95 237 -75
rect 249 -95 253 -75
rect 257 -95 261 -75
rect 6 -132 10 -112
rect 17 -132 21 -112
rect 28 -132 32 -112
rect 44 -132 48 -112
rect 52 -132 56 -112
rect 6 -223 10 -203
rect 17 -223 21 -203
rect 28 -223 32 -203
rect 44 -223 48 -203
rect 52 -223 56 -203
rect 68 -223 72 -203
rect 79 -223 83 -203
rect 90 -223 94 -203
rect 106 -223 110 -203
rect 114 -223 118 -203
rect 130 -223 134 -203
rect 141 -223 145 -203
rect 152 -223 156 -203
rect 168 -223 172 -203
rect 176 -223 180 -203
rect 6 -320 10 -300
rect 17 -320 21 -300
rect 28 -320 32 -300
rect 44 -320 48 -300
rect 52 -320 56 -300
rect 68 -320 72 -300
rect 79 -320 83 -300
rect 90 -320 94 -300
rect 106 -320 110 -300
rect 114 -320 118 -300
rect 236 -307 240 -287
rect 258 -307 262 -287
rect 274 -307 278 -287
rect 282 -307 286 -287
rect 298 -307 302 -287
rect 320 -307 324 -287
rect 336 -307 340 -287
rect 344 -307 348 -287
rect 360 -307 364 -287
rect 382 -307 386 -287
rect 398 -307 402 -287
rect 406 -307 410 -287
rect 6 -405 10 -385
rect 17 -405 21 -385
rect 28 -405 32 -385
rect 44 -405 48 -385
rect 52 -405 56 -385
rect 6 -517 10 -497
rect 17 -517 21 -497
rect 28 -517 32 -497
rect 44 -517 48 -497
rect 52 -517 56 -497
rect 68 -517 72 -497
rect 79 -517 83 -497
rect 90 -517 94 -497
rect 106 -517 110 -497
rect 114 -517 118 -497
rect 130 -517 134 -497
rect 141 -517 145 -497
rect 152 -517 156 -497
rect 168 -517 172 -497
rect 176 -517 180 -497
rect 192 -517 196 -497
rect 203 -517 207 -497
rect 214 -517 218 -497
rect 230 -517 234 -497
rect 238 -517 242 -497
rect 6 -617 10 -597
rect 17 -617 21 -597
rect 28 -617 32 -597
rect 44 -617 48 -597
rect 52 -617 56 -597
rect 68 -617 72 -597
rect 79 -617 83 -597
rect 90 -617 94 -597
rect 106 -617 110 -597
rect 114 -617 118 -597
rect 130 -617 134 -597
rect 141 -617 145 -597
rect 152 -617 156 -597
rect 168 -617 172 -597
rect 176 -617 180 -597
rect 6 -717 10 -697
rect 17 -717 21 -697
rect 28 -717 32 -697
rect 44 -717 48 -697
rect 52 -717 56 -697
rect 68 -717 72 -697
rect 79 -717 83 -697
rect 90 -717 94 -697
rect 106 -717 110 -697
rect 114 -717 118 -697
rect 314 -699 318 -679
rect 336 -699 340 -679
rect 352 -699 356 -679
rect 360 -699 364 -679
rect 376 -699 380 -679
rect 398 -699 402 -679
rect 414 -699 418 -679
rect 422 -699 426 -679
rect 438 -699 442 -679
rect 460 -699 464 -679
rect 476 -699 480 -679
rect 484 -699 488 -679
rect 500 -699 504 -679
rect 522 -699 526 -679
rect 538 -699 542 -679
rect 546 -699 550 -679
rect 6 -817 10 -797
rect 17 -817 21 -797
rect 28 -817 32 -797
rect 44 -817 48 -797
rect 52 -817 56 -797
<< psubstratepcontact >>
rect 48 0 52 4
rect 110 -6 114 -2
rect 48 -89 52 -85
rect 110 -89 114 -85
rect 191 -141 195 -137
rect 253 -141 257 -137
rect 48 -172 52 -168
rect 48 -263 52 -259
rect 110 -263 114 -259
rect 172 -263 176 -259
rect 278 -353 282 -349
rect 340 -353 344 -349
rect 402 -353 406 -349
rect 48 -360 52 -356
rect 110 -360 114 -356
rect 48 -445 52 -441
rect 48 -557 52 -553
rect 110 -557 114 -553
rect 172 -557 176 -553
rect 234 -557 238 -553
rect 48 -657 52 -653
rect 110 -657 114 -653
rect 172 -657 176 -653
rect 356 -745 360 -741
rect 418 -745 422 -741
rect 480 -745 484 -741
rect 542 -745 546 -741
rect 48 -757 52 -753
rect 110 -757 114 -753
rect 48 -857 52 -853
<< nsubstratencontact >>
rect 48 64 52 68
rect 110 64 114 68
rect 48 -25 52 -21
rect 110 -25 114 -21
rect 191 -71 195 -67
rect 253 -71 257 -67
rect 48 -108 52 -104
rect 48 -199 52 -195
rect 110 -199 114 -195
rect 172 -199 176 -195
rect 278 -283 282 -279
rect 340 -283 344 -279
rect 402 -283 406 -279
rect 48 -296 52 -292
rect 110 -296 114 -292
rect 48 -381 52 -377
rect 48 -493 52 -489
rect 110 -493 114 -489
rect 172 -493 176 -489
rect 234 -493 238 -489
rect 48 -593 52 -589
rect 110 -593 114 -589
rect 172 -593 176 -589
rect 356 -675 360 -671
rect 418 -675 422 -671
rect 480 -675 484 -671
rect 542 -675 546 -671
rect 48 -693 52 -689
rect 110 -693 114 -689
rect 48 -793 52 -789
<< polysilicon >>
rect 11 60 13 63
rect 25 60 27 63
rect 49 60 51 63
rect 73 60 75 63
rect 87 60 89 63
rect 111 60 113 63
rect 11 18 13 40
rect 25 18 27 40
rect 49 18 51 40
rect 73 12 75 40
rect 87 12 89 40
rect 111 12 113 40
rect 11 5 13 8
rect 25 5 27 8
rect 49 5 51 8
rect 73 -1 75 2
rect 87 -1 89 2
rect 111 -1 113 2
rect 11 -29 13 -26
rect 25 -29 27 -26
rect 49 -29 51 -26
rect 73 -29 75 -26
rect 87 -29 89 -26
rect 111 -29 113 -26
rect 11 -71 13 -49
rect 25 -71 27 -49
rect 49 -71 51 -49
rect 73 -71 75 -49
rect 87 -71 89 -49
rect 111 -71 113 -49
rect 154 -75 156 -72
rect 168 -75 170 -72
rect 192 -75 194 -72
rect 216 -75 218 -72
rect 230 -75 232 -72
rect 254 -75 256 -72
rect 11 -84 13 -81
rect 25 -84 27 -81
rect 49 -84 51 -81
rect 73 -84 75 -81
rect 87 -84 89 -81
rect 111 -84 113 -81
rect 11 -112 13 -109
rect 25 -112 27 -109
rect 49 -112 51 -109
rect 154 -123 156 -95
rect 168 -123 170 -95
rect 192 -123 194 -95
rect 216 -123 218 -95
rect 230 -123 232 -95
rect 254 -123 256 -95
rect 11 -154 13 -132
rect 25 -154 27 -132
rect 49 -154 51 -132
rect 154 -136 156 -133
rect 168 -136 170 -133
rect 192 -136 194 -133
rect 216 -136 218 -133
rect 230 -136 232 -133
rect 254 -136 256 -133
rect 11 -167 13 -164
rect 25 -167 27 -164
rect 49 -167 51 -164
rect 11 -203 13 -200
rect 25 -203 27 -200
rect 49 -203 51 -200
rect 73 -203 75 -200
rect 87 -203 89 -200
rect 111 -203 113 -200
rect 135 -203 137 -200
rect 149 -203 151 -200
rect 173 -203 175 -200
rect 11 -245 13 -223
rect 25 -245 27 -223
rect 49 -245 51 -223
rect 73 -245 75 -223
rect 87 -245 89 -223
rect 111 -245 113 -223
rect 135 -245 137 -223
rect 149 -245 151 -223
rect 173 -245 175 -223
rect 11 -258 13 -255
rect 25 -258 27 -255
rect 49 -258 51 -255
rect 73 -258 75 -255
rect 87 -258 89 -255
rect 111 -258 113 -255
rect 135 -258 137 -255
rect 149 -258 151 -255
rect 173 -258 175 -255
rect 241 -287 243 -284
rect 255 -287 257 -284
rect 279 -287 281 -284
rect 303 -287 305 -284
rect 317 -287 319 -284
rect 341 -287 343 -284
rect 365 -287 367 -284
rect 379 -287 381 -284
rect 403 -287 405 -284
rect 11 -300 13 -297
rect 25 -300 27 -297
rect 49 -300 51 -297
rect 73 -300 75 -297
rect 87 -300 89 -297
rect 111 -300 113 -297
rect 11 -342 13 -320
rect 25 -342 27 -320
rect 49 -342 51 -320
rect 73 -342 75 -320
rect 87 -342 89 -320
rect 111 -342 113 -320
rect 241 -335 243 -307
rect 255 -335 257 -307
rect 279 -335 281 -307
rect 303 -335 305 -307
rect 317 -335 319 -307
rect 341 -335 343 -307
rect 365 -335 367 -307
rect 379 -335 381 -307
rect 403 -335 405 -307
rect 241 -348 243 -345
rect 255 -348 257 -345
rect 279 -348 281 -345
rect 303 -348 305 -345
rect 317 -348 319 -345
rect 341 -348 343 -345
rect 365 -348 367 -345
rect 379 -348 381 -345
rect 403 -348 405 -345
rect 11 -355 13 -352
rect 25 -355 27 -352
rect 49 -355 51 -352
rect 73 -355 75 -352
rect 87 -355 89 -352
rect 111 -355 113 -352
rect 11 -385 13 -382
rect 25 -385 27 -382
rect 49 -385 51 -382
rect 11 -427 13 -405
rect 25 -427 27 -405
rect 49 -427 51 -405
rect 11 -440 13 -437
rect 25 -440 27 -437
rect 49 -440 51 -437
rect 11 -497 13 -494
rect 25 -497 27 -494
rect 49 -497 51 -494
rect 73 -497 75 -494
rect 87 -497 89 -494
rect 111 -497 113 -494
rect 135 -497 137 -494
rect 149 -497 151 -494
rect 173 -497 175 -494
rect 197 -497 199 -494
rect 211 -497 213 -494
rect 235 -497 237 -494
rect 11 -539 13 -517
rect 25 -539 27 -517
rect 49 -539 51 -517
rect 73 -539 75 -517
rect 87 -539 89 -517
rect 111 -539 113 -517
rect 135 -539 137 -517
rect 149 -539 151 -517
rect 173 -539 175 -517
rect 197 -539 199 -517
rect 211 -539 213 -517
rect 235 -539 237 -517
rect 11 -552 13 -549
rect 25 -552 27 -549
rect 49 -552 51 -549
rect 73 -552 75 -549
rect 87 -552 89 -549
rect 111 -552 113 -549
rect 135 -552 137 -549
rect 149 -552 151 -549
rect 173 -552 175 -549
rect 197 -552 199 -549
rect 211 -552 213 -549
rect 235 -552 237 -549
rect 11 -597 13 -594
rect 25 -597 27 -594
rect 49 -597 51 -594
rect 73 -597 75 -594
rect 87 -597 89 -594
rect 111 -597 113 -594
rect 135 -597 137 -594
rect 149 -597 151 -594
rect 173 -597 175 -594
rect 11 -639 13 -617
rect 25 -639 27 -617
rect 49 -639 51 -617
rect 73 -639 75 -617
rect 87 -639 89 -617
rect 111 -639 113 -617
rect 135 -639 137 -617
rect 149 -639 151 -617
rect 173 -639 175 -617
rect 11 -652 13 -649
rect 25 -652 27 -649
rect 49 -652 51 -649
rect 73 -652 75 -649
rect 87 -652 89 -649
rect 111 -652 113 -649
rect 135 -652 137 -649
rect 149 -652 151 -649
rect 173 -652 175 -649
rect 319 -679 321 -676
rect 333 -679 335 -676
rect 357 -679 359 -676
rect 381 -679 383 -676
rect 395 -679 397 -676
rect 419 -679 421 -676
rect 443 -679 445 -676
rect 457 -679 459 -676
rect 481 -679 483 -676
rect 505 -679 507 -676
rect 519 -679 521 -676
rect 543 -679 545 -676
rect 11 -697 13 -694
rect 25 -697 27 -694
rect 49 -697 51 -694
rect 73 -697 75 -694
rect 87 -697 89 -694
rect 111 -697 113 -694
rect 11 -739 13 -717
rect 25 -739 27 -717
rect 49 -739 51 -717
rect 73 -739 75 -717
rect 87 -739 89 -717
rect 111 -739 113 -717
rect 319 -727 321 -699
rect 333 -727 335 -699
rect 357 -727 359 -699
rect 381 -727 383 -699
rect 395 -727 397 -699
rect 419 -727 421 -699
rect 443 -727 445 -699
rect 457 -727 459 -699
rect 481 -727 483 -699
rect 505 -727 507 -699
rect 519 -727 521 -699
rect 543 -727 545 -699
rect 319 -740 321 -737
rect 333 -740 335 -737
rect 357 -740 359 -737
rect 381 -740 383 -737
rect 395 -740 397 -737
rect 419 -740 421 -737
rect 443 -740 445 -737
rect 457 -740 459 -737
rect 481 -740 483 -737
rect 505 -740 507 -737
rect 519 -740 521 -737
rect 543 -740 545 -737
rect 11 -752 13 -749
rect 25 -752 27 -749
rect 49 -752 51 -749
rect 73 -752 75 -749
rect 87 -752 89 -749
rect 111 -752 113 -749
rect 11 -797 13 -794
rect 25 -797 27 -794
rect 49 -797 51 -794
rect 11 -839 13 -817
rect 25 -839 27 -817
rect 49 -839 51 -817
rect 11 -852 13 -849
rect 25 -852 27 -849
rect 49 -852 51 -849
<< polycontact >>
rect 7 29 11 33
rect 21 22 25 26
rect 45 29 49 33
rect 69 29 73 33
rect 83 22 87 26
rect 107 29 111 33
rect 7 -60 11 -56
rect 21 -67 25 -63
rect 45 -60 49 -56
rect 69 -60 73 -56
rect 83 -67 87 -63
rect 107 -60 111 -56
rect 150 -106 154 -102
rect 164 -113 168 -109
rect 188 -106 192 -102
rect 212 -106 216 -102
rect 226 -113 230 -109
rect 250 -106 254 -102
rect 7 -143 11 -139
rect 21 -150 25 -146
rect 45 -143 49 -139
rect 7 -234 11 -230
rect 21 -241 25 -237
rect 45 -234 49 -230
rect 69 -234 73 -230
rect 83 -241 87 -237
rect 107 -234 111 -230
rect 131 -234 135 -230
rect 145 -241 149 -237
rect 169 -234 173 -230
rect 237 -318 241 -314
rect 7 -331 11 -327
rect 21 -338 25 -334
rect 45 -331 49 -327
rect 69 -331 73 -327
rect 83 -338 87 -334
rect 107 -331 111 -327
rect 251 -325 255 -321
rect 275 -318 279 -314
rect 299 -318 303 -314
rect 313 -325 317 -321
rect 337 -318 341 -314
rect 361 -318 365 -314
rect 375 -325 379 -321
rect 399 -318 403 -314
rect 7 -416 11 -412
rect 21 -423 25 -419
rect 45 -416 49 -412
rect 7 -528 11 -524
rect 21 -535 25 -531
rect 45 -528 49 -524
rect 69 -528 73 -524
rect 83 -535 87 -531
rect 107 -528 111 -524
rect 131 -528 135 -524
rect 145 -535 149 -531
rect 169 -528 173 -524
rect 193 -528 197 -524
rect 207 -535 211 -531
rect 231 -528 235 -524
rect 7 -628 11 -624
rect 21 -635 25 -631
rect 45 -628 49 -624
rect 69 -628 73 -624
rect 83 -635 87 -631
rect 107 -628 111 -624
rect 131 -628 135 -624
rect 145 -635 149 -631
rect 169 -628 173 -624
rect 315 -710 319 -706
rect 7 -728 11 -724
rect 21 -735 25 -731
rect 45 -728 49 -724
rect 69 -728 73 -724
rect 83 -735 87 -731
rect 107 -728 111 -724
rect 329 -717 333 -713
rect 353 -710 357 -706
rect 377 -710 381 -706
rect 391 -717 395 -713
rect 415 -710 419 -706
rect 439 -710 443 -706
rect 453 -717 457 -713
rect 477 -710 481 -706
rect 501 -710 505 -706
rect 515 -717 519 -713
rect 539 -710 543 -706
rect 7 -828 11 -824
rect 21 -835 25 -831
rect 45 -828 49 -824
<< metal1 >>
rect 6 68 119 70
rect 6 64 48 68
rect 52 64 110 68
rect 114 64 119 68
rect 6 60 10 64
rect 28 60 32 64
rect 44 60 48 64
rect 68 60 72 64
rect 106 60 110 64
rect 17 33 21 40
rect 52 33 56 40
rect 90 33 94 40
rect 114 33 118 40
rect -15 29 7 33
rect 17 29 45 33
rect 52 29 69 33
rect 90 29 107 33
rect 114 29 124 33
rect -30 21 -25 26
rect -15 -56 -11 29
rect 4 22 21 26
rect 28 18 32 29
rect 52 18 56 29
rect 65 22 83 26
rect 90 19 94 29
rect 68 15 94 19
rect 68 12 72 15
rect 90 12 94 15
rect 114 12 118 29
rect 6 4 10 8
rect 44 4 48 8
rect 6 0 16 4
rect 21 0 48 4
rect 52 0 60 4
rect 56 -2 60 0
rect 79 -2 83 2
rect 106 -2 110 2
rect 56 -6 110 -2
rect 114 -6 141 -2
rect 0 -15 60 -10
rect 6 -21 119 -19
rect 6 -25 48 -21
rect 52 -25 110 -21
rect 114 -25 119 -21
rect 6 -29 10 -25
rect 28 -29 32 -25
rect 44 -29 48 -25
rect 68 -29 72 -25
rect 90 -29 94 -25
rect 106 -29 110 -25
rect 17 -56 21 -49
rect 52 -56 56 -49
rect 79 -56 83 -49
rect 114 -56 118 -49
rect -15 -60 7 -56
rect 17 -60 45 -56
rect 52 -60 69 -56
rect 79 -60 107 -56
rect 114 -60 135 -56
rect -15 -230 -11 -60
rect 0 -64 21 -63
rect 3 -67 21 -64
rect 28 -71 32 -60
rect 52 -71 56 -60
rect 66 -67 83 -63
rect 90 -71 94 -60
rect 114 -71 118 -60
rect 6 -85 10 -81
rect 6 -89 16 -85
rect 44 -85 48 -81
rect 68 -85 72 -81
rect 106 -85 110 -81
rect 21 -89 48 -85
rect 52 -89 110 -85
rect 114 -89 124 -85
rect -3 -98 61 -93
rect -3 -139 2 -98
rect 131 -102 135 -60
rect 143 -71 153 -65
rect 159 -67 267 -65
rect 159 -71 191 -67
rect 195 -71 253 -67
rect 257 -71 267 -67
rect 149 -75 153 -71
rect 187 -75 191 -71
rect 211 -75 215 -71
rect 249 -75 253 -71
rect 171 -102 175 -95
rect 195 -102 199 -95
rect 233 -102 237 -95
rect 257 -102 261 -95
rect 6 -104 56 -102
rect 6 -108 48 -104
rect 52 -108 56 -104
rect 131 -106 150 -102
rect 171 -106 188 -102
rect 195 -106 212 -102
rect 233 -106 250 -102
rect 257 -106 267 -102
rect 6 -112 10 -108
rect 28 -112 32 -108
rect 44 -112 48 -108
rect 17 -139 21 -132
rect 52 -139 56 -132
rect 131 -113 164 -109
rect 131 -139 135 -113
rect 171 -116 175 -106
rect 149 -120 175 -116
rect 149 -123 153 -120
rect 171 -123 175 -120
rect 195 -123 199 -106
rect 208 -113 226 -109
rect 233 -116 237 -106
rect 211 -120 237 -116
rect 211 -123 215 -120
rect 233 -123 237 -120
rect 257 -123 261 -106
rect -3 -143 7 -139
rect 17 -143 45 -139
rect 52 -143 135 -139
rect 160 -137 164 -133
rect 187 -137 191 -133
rect 222 -137 226 -133
rect 249 -137 253 -133
rect 160 -141 191 -137
rect 195 -141 253 -137
rect 257 -141 262 -137
rect 0 -150 21 -146
rect 28 -154 32 -143
rect 52 -154 56 -143
rect 171 -150 203 -145
rect 6 -168 10 -164
rect 6 -172 16 -168
rect 44 -168 48 -164
rect 21 -172 48 -168
rect 6 -195 128 -193
rect 6 -199 48 -195
rect 52 -199 110 -195
rect 114 -199 128 -195
rect 134 -195 186 -193
rect 134 -199 172 -195
rect 176 -199 186 -195
rect 6 -203 10 -199
rect 28 -203 32 -199
rect 44 -203 48 -199
rect 68 -203 72 -199
rect 90 -203 94 -199
rect 106 -203 110 -199
rect 130 -203 134 -199
rect 152 -203 156 -199
rect 168 -203 172 -199
rect 17 -230 21 -223
rect 52 -230 56 -223
rect 79 -230 83 -223
rect 114 -230 118 -223
rect 141 -230 145 -223
rect 176 -230 180 -223
rect -15 -234 7 -230
rect 17 -234 45 -230
rect 52 -234 69 -230
rect 79 -234 107 -230
rect 114 -234 131 -230
rect 141 -234 169 -230
rect 176 -234 209 -230
rect -15 -524 -11 -234
rect -2 -238 21 -237
rect 2 -241 21 -238
rect 28 -245 32 -234
rect 52 -245 56 -234
rect 65 -241 83 -237
rect 90 -245 94 -234
rect 114 -245 118 -234
rect 128 -241 145 -237
rect 152 -245 156 -234
rect 176 -245 180 -234
rect 6 -259 10 -255
rect 6 -263 16 -259
rect 44 -259 48 -255
rect 68 -259 72 -255
rect 106 -259 110 -255
rect 130 -259 134 -255
rect 168 -259 172 -255
rect 21 -263 48 -259
rect 52 -263 110 -259
rect 114 -263 172 -259
rect 176 -263 186 -259
rect -7 -272 60 -267
rect 114 -272 123 -267
rect -7 -327 -2 -272
rect 6 -292 119 -290
rect 6 -296 48 -292
rect 52 -296 110 -292
rect 114 -296 119 -292
rect 6 -300 10 -296
rect 28 -300 32 -296
rect 44 -300 48 -296
rect 68 -300 72 -296
rect 90 -300 94 -296
rect 106 -300 110 -296
rect 205 -314 209 -234
rect 230 -283 231 -277
rect 237 -279 416 -277
rect 237 -283 278 -279
rect 282 -283 340 -279
rect 344 -283 402 -279
rect 406 -283 416 -279
rect 236 -287 240 -283
rect 274 -287 278 -283
rect 298 -287 302 -283
rect 336 -287 340 -283
rect 360 -287 364 -283
rect 398 -287 402 -283
rect 258 -314 262 -307
rect 282 -314 286 -307
rect 320 -314 324 -307
rect 344 -314 348 -307
rect 382 -314 386 -307
rect 406 -314 410 -307
rect 205 -318 237 -314
rect 258 -318 275 -314
rect 282 -318 299 -314
rect 320 -318 337 -314
rect 344 -318 361 -314
rect 382 -318 399 -314
rect 406 -318 416 -314
rect 17 -327 21 -320
rect 52 -327 56 -320
rect 79 -327 83 -320
rect 114 -327 118 -320
rect 205 -325 251 -321
rect 205 -327 209 -325
rect -7 -331 7 -327
rect 17 -331 45 -327
rect 52 -331 69 -327
rect 79 -331 107 -327
rect 114 -331 209 -327
rect 258 -328 262 -318
rect 0 -338 21 -334
rect 28 -342 32 -331
rect 52 -342 56 -331
rect 65 -338 83 -334
rect 90 -342 94 -331
rect 114 -342 118 -331
rect 236 -332 262 -328
rect 236 -335 240 -332
rect 258 -335 262 -332
rect 282 -335 286 -318
rect 295 -325 313 -321
rect 320 -328 324 -318
rect 298 -332 324 -328
rect 298 -335 302 -332
rect 320 -335 324 -332
rect 344 -335 348 -318
rect 357 -325 375 -321
rect 382 -328 386 -318
rect 360 -332 386 -328
rect 360 -335 364 -332
rect 382 -335 386 -332
rect 406 -335 410 -318
rect 247 -349 251 -345
rect 274 -349 278 -345
rect 309 -349 313 -345
rect 336 -349 340 -345
rect 371 -349 375 -345
rect 398 -349 402 -345
rect 6 -356 10 -352
rect 6 -360 16 -356
rect 44 -356 48 -352
rect 68 -356 72 -352
rect 106 -356 110 -352
rect 233 -353 278 -349
rect 282 -353 340 -349
rect 344 -353 402 -349
rect 406 -353 411 -349
rect 21 -360 48 -356
rect 52 -360 110 -356
rect 114 -360 124 -356
rect 239 -362 290 -357
rect 345 -362 352 -357
rect 52 -369 60 -364
rect 6 -377 57 -375
rect 6 -381 48 -377
rect 52 -381 57 -377
rect 6 -385 10 -381
rect 28 -385 32 -381
rect 44 -385 48 -381
rect 17 -412 21 -405
rect 52 -412 56 -405
rect 239 -412 243 -362
rect 0 -416 7 -412
rect 17 -416 45 -412
rect 52 -416 243 -412
rect 0 -423 21 -419
rect 28 -427 32 -416
rect 52 -427 56 -416
rect 6 -441 10 -437
rect 6 -445 16 -441
rect 44 -441 48 -437
rect 21 -445 48 -441
rect 52 -445 60 -441
rect 6 -489 193 -487
rect 6 -493 48 -489
rect 52 -493 110 -489
rect 114 -493 172 -489
rect 176 -493 193 -489
rect 199 -489 248 -487
rect 199 -493 234 -489
rect 238 -493 248 -489
rect 6 -497 10 -493
rect 28 -497 32 -493
rect 44 -497 48 -493
rect 68 -497 72 -493
rect 90 -497 94 -493
rect 106 -497 110 -493
rect 130 -497 134 -493
rect 152 -497 156 -493
rect 168 -497 172 -493
rect 192 -497 196 -493
rect 214 -497 218 -493
rect 230 -497 234 -493
rect 17 -524 21 -517
rect 52 -524 56 -517
rect 79 -524 83 -517
rect 114 -524 118 -517
rect 141 -524 145 -517
rect 176 -524 180 -517
rect 203 -524 207 -517
rect 238 -524 242 -517
rect -15 -528 7 -524
rect 17 -528 45 -524
rect 52 -528 69 -524
rect 79 -528 107 -524
rect 114 -528 131 -524
rect 141 -528 169 -524
rect 176 -528 193 -524
rect 203 -528 231 -524
rect 238 -528 264 -524
rect 3 -535 21 -531
rect 28 -539 32 -528
rect 52 -539 56 -528
rect 66 -535 83 -531
rect 90 -539 94 -528
rect 114 -539 118 -528
rect 127 -535 145 -531
rect 152 -539 156 -528
rect 176 -539 180 -528
rect 189 -535 207 -531
rect 214 -539 218 -528
rect 238 -539 242 -528
rect 6 -553 10 -549
rect 6 -557 16 -553
rect 44 -553 48 -549
rect 68 -553 72 -549
rect 106 -553 110 -549
rect 130 -553 134 -549
rect 168 -553 172 -549
rect 192 -553 196 -549
rect 230 -553 234 -549
rect 21 -557 48 -553
rect 52 -557 110 -553
rect 114 -557 172 -553
rect 176 -557 234 -553
rect 238 -557 248 -553
rect 56 -566 61 -561
rect 116 -566 122 -561
rect 178 -566 184 -561
rect 6 -589 181 -587
rect 6 -593 48 -589
rect 52 -593 110 -589
rect 114 -593 172 -589
rect 176 -593 181 -589
rect 6 -597 10 -593
rect 28 -597 32 -593
rect 44 -597 48 -593
rect 68 -597 72 -593
rect 90 -597 94 -593
rect 106 -597 110 -593
rect 130 -597 134 -593
rect 152 -597 156 -593
rect 168 -597 172 -593
rect 17 -624 21 -617
rect 52 -624 56 -617
rect 79 -624 83 -617
rect 114 -624 118 -617
rect 141 -624 145 -617
rect 176 -624 180 -617
rect 0 -628 7 -624
rect 17 -628 45 -624
rect 52 -628 69 -624
rect 79 -628 107 -624
rect 114 -628 131 -624
rect 141 -628 169 -624
rect 176 -628 233 -624
rect 0 -635 21 -631
rect 28 -639 32 -628
rect 52 -639 56 -628
rect 66 -635 83 -631
rect 90 -639 94 -628
rect 114 -639 118 -628
rect 127 -635 145 -631
rect 152 -639 156 -628
rect 176 -639 180 -628
rect 6 -653 10 -649
rect 6 -657 16 -653
rect 44 -653 48 -649
rect 68 -653 72 -649
rect 106 -653 110 -649
rect 130 -653 134 -649
rect 168 -653 172 -649
rect 21 -657 48 -653
rect 52 -657 110 -653
rect 114 -657 172 -653
rect 176 -657 186 -653
rect 56 -666 61 -661
rect 116 -666 122 -661
rect 6 -689 119 -687
rect 6 -693 48 -689
rect 52 -693 110 -689
rect 114 -693 119 -689
rect 6 -697 10 -693
rect 28 -697 32 -693
rect 44 -697 48 -693
rect 68 -697 72 -693
rect 90 -697 94 -693
rect 106 -697 110 -693
rect 229 -713 233 -628
rect 260 -706 264 -528
rect 308 -675 328 -669
rect 334 -671 556 -669
rect 334 -675 356 -671
rect 360 -675 418 -671
rect 422 -675 480 -671
rect 484 -675 542 -671
rect 546 -675 556 -671
rect 314 -679 318 -675
rect 352 -679 356 -675
rect 376 -679 380 -675
rect 414 -679 418 -675
rect 438 -679 442 -675
rect 476 -679 480 -675
rect 500 -679 504 -675
rect 538 -679 542 -675
rect 336 -706 340 -699
rect 360 -706 364 -699
rect 398 -706 402 -699
rect 422 -706 426 -699
rect 460 -706 464 -699
rect 484 -706 488 -699
rect 522 -706 526 -699
rect 546 -706 550 -699
rect 260 -710 315 -706
rect 336 -710 353 -706
rect 360 -710 377 -706
rect 398 -710 415 -706
rect 422 -710 439 -706
rect 460 -710 477 -706
rect 484 -710 501 -706
rect 522 -710 539 -706
rect 546 -710 556 -706
rect 229 -717 329 -713
rect 17 -724 21 -717
rect 52 -724 56 -717
rect 79 -724 83 -717
rect 114 -724 118 -717
rect 336 -720 340 -710
rect 314 -724 340 -720
rect 0 -728 7 -724
rect 17 -728 45 -724
rect 52 -728 69 -724
rect 79 -728 107 -724
rect 114 -728 233 -724
rect 0 -735 21 -731
rect 28 -739 32 -728
rect 52 -739 56 -728
rect 66 -735 83 -731
rect 90 -739 94 -728
rect 114 -739 118 -728
rect 229 -749 233 -728
rect 314 -727 318 -724
rect 336 -727 340 -724
rect 360 -727 364 -710
rect 373 -717 391 -713
rect 398 -720 402 -710
rect 376 -724 402 -720
rect 376 -727 380 -724
rect 398 -727 402 -724
rect 422 -727 426 -710
rect 435 -717 453 -713
rect 460 -720 464 -710
rect 438 -724 464 -720
rect 438 -727 442 -724
rect 460 -727 464 -724
rect 484 -727 488 -710
rect 497 -717 515 -713
rect 522 -720 526 -710
rect 500 -724 526 -720
rect 500 -727 504 -724
rect 522 -727 526 -724
rect 546 -727 550 -710
rect 325 -741 329 -737
rect 352 -741 356 -737
rect 387 -741 391 -737
rect 414 -741 418 -737
rect 449 -741 453 -737
rect 476 -741 480 -737
rect 511 -741 515 -737
rect 538 -741 542 -737
rect 311 -745 356 -741
rect 360 -745 418 -741
rect 422 -745 480 -741
rect 484 -745 542 -741
rect 546 -745 551 -741
rect 6 -753 10 -749
rect 6 -757 16 -753
rect 44 -753 48 -749
rect 68 -753 72 -749
rect 106 -753 110 -749
rect 21 -757 48 -753
rect 52 -757 110 -753
rect 114 -757 124 -753
rect 229 -754 368 -749
rect 486 -754 492 -749
rect 56 -766 61 -761
rect 6 -789 57 -787
rect 6 -793 48 -789
rect 52 -793 57 -789
rect 6 -797 10 -793
rect 28 -797 32 -793
rect 44 -797 48 -793
rect 17 -824 21 -817
rect 52 -824 56 -817
rect 430 -824 435 -754
rect 0 -828 7 -824
rect 17 -828 45 -824
rect 52 -828 435 -824
rect 0 -835 21 -831
rect 28 -839 32 -828
rect 52 -839 56 -828
rect 6 -853 10 -849
rect 6 -857 16 -853
rect 44 -853 48 -849
rect 21 -857 48 -853
rect 52 -857 62 -853
<< m2contact >>
rect 119 64 124 70
rect -25 21 -20 26
rect -1 21 4 26
rect 60 21 65 26
rect 16 -1 21 4
rect 141 -6 146 -1
rect 60 -15 65 -10
rect 119 -25 124 -19
rect -2 -69 3 -64
rect 61 -68 66 -63
rect 16 -89 21 -84
rect 61 -98 66 -93
rect 153 -71 159 -65
rect 56 -108 62 -102
rect 203 -114 208 -109
rect 262 -141 267 -136
rect 203 -150 208 -145
rect 16 -172 21 -167
rect 128 -199 134 -193
rect -3 -243 2 -238
rect 60 -242 65 -237
rect 123 -242 128 -237
rect 16 -263 21 -258
rect 60 -272 65 -267
rect 123 -272 128 -267
rect 119 -296 124 -290
rect 231 -283 237 -277
rect 60 -339 65 -334
rect 290 -326 295 -321
rect 352 -326 357 -321
rect 16 -360 21 -355
rect 411 -353 416 -348
rect 290 -362 295 -357
rect 352 -362 357 -357
rect 60 -369 65 -364
rect 57 -381 62 -375
rect 16 -445 21 -440
rect 193 -493 199 -487
rect -2 -537 3 -531
rect 61 -536 66 -531
rect 122 -536 127 -531
rect 184 -536 189 -531
rect 16 -557 21 -552
rect 61 -566 66 -561
rect 122 -566 127 -561
rect 184 -566 189 -561
rect 181 -593 186 -587
rect 61 -636 66 -631
rect 122 -636 127 -631
rect 16 -657 21 -652
rect 61 -666 66 -661
rect 122 -666 127 -661
rect 119 -693 124 -687
rect 328 -675 334 -669
rect 61 -736 66 -731
rect 368 -718 373 -713
rect 430 -718 435 -713
rect 492 -718 497 -713
rect 551 -745 556 -740
rect 16 -757 21 -752
rect 368 -754 373 -749
rect 430 -754 435 -749
rect 492 -754 497 -749
rect 61 -766 66 -761
rect 57 -793 62 -787
rect 16 -857 21 -852
<< metal2 >>
rect 124 64 134 70
rect -20 21 -1 26
rect -15 -64 -10 21
rect -15 -69 -2 -64
rect -15 -238 -10 -69
rect 16 -84 21 -1
rect 60 -10 65 21
rect 128 -19 134 64
rect 146 -6 293 -1
rect 124 -25 159 -19
rect 16 -167 21 -89
rect 61 -93 66 -68
rect 128 -102 134 -25
rect 153 -65 159 -25
rect 62 -108 134 -102
rect -15 -243 -3 -238
rect -15 -532 -10 -243
rect 16 -258 21 -172
rect 128 -176 134 -108
rect 203 -145 208 -114
rect 288 -136 293 -6
rect 267 -141 454 -136
rect 128 -182 237 -176
rect 128 -193 134 -182
rect 16 -355 21 -263
rect 60 -267 65 -242
rect 123 -267 128 -242
rect 231 -270 237 -182
rect 193 -276 237 -270
rect 193 -290 199 -276
rect 231 -277 237 -276
rect 124 -296 199 -290
rect 16 -440 21 -360
rect 60 -364 65 -339
rect 193 -375 199 -296
rect 290 -357 295 -326
rect 352 -357 357 -326
rect 449 -346 454 -141
rect 449 -348 615 -346
rect 416 -351 615 -348
rect 416 -353 454 -351
rect 62 -381 199 -375
rect -15 -537 -2 -532
rect 16 -552 21 -445
rect 193 -474 199 -381
rect 193 -480 334 -474
rect 193 -487 199 -480
rect 16 -652 21 -557
rect 61 -561 66 -536
rect 122 -561 127 -536
rect 184 -561 189 -536
rect 328 -587 334 -480
rect 186 -593 334 -587
rect 16 -752 21 -657
rect 61 -661 66 -636
rect 122 -661 127 -636
rect 209 -687 215 -593
rect 328 -669 334 -593
rect 124 -693 215 -687
rect 16 -852 21 -757
rect 61 -761 66 -736
rect 138 -787 144 -693
rect 368 -749 373 -718
rect 430 -749 435 -718
rect 492 -749 497 -718
rect 610 -740 615 -351
rect 556 -745 615 -740
rect 62 -793 144 -787
<< labels >>
rlabel metal1 122 31 122 31 1 C1
rlabel metal1 266 -104 266 -104 7 C2
rlabel metal1 415 -316 415 -316 1 C3
rlabel metal1 554 -708 554 -708 7 Cout
rlabel metal1 35 -855 35 -855 1 gnd
rlabel metal1 61 67 61 67 5 vdd
rlabel metal1 -13 31 -13 31 3 Cin
rlabel metal1 -29 23 -29 23 3 P0
rlabel metal1 3 -13 3 -13 1 G0
rlabel metal1 0 -96 0 -96 1 P1
rlabel metal1 2 -148 2 -148 1 G0
rlabel metal1 174 -148 174 -148 1 G1
rlabel metal1 116 -270 116 -270 1 P2
rlabel metal1 52 -270 52 -270 1 P1
rlabel metal1 3 -336 3 -336 1 P2
rlabel metal1 54 -367 54 -367 1 G0
rlabel metal1 2 -414 2 -414 1 P2
rlabel metal1 2 -421 2 -421 1 G1
rlabel metal1 347 -360 347 -360 1 G2
rlabel metal1 58 -564 58 -564 1 P1
rlabel metal1 2 -626 2 -626 1 P1
rlabel metal1 118 -563 118 -563 1 P2
rlabel metal1 2 -633 2 -633 1 P2
rlabel metal1 179 -564 179 -564 1 P3
rlabel metal1 57 -664 57 -664 1 P3
rlabel metal1 117 -664 117 -664 1 G0
rlabel metal1 2 -726 2 -726 1 P3
rlabel metal1 2 -733 2 -733 1 P2
rlabel metal1 58 -764 58 -764 1 G1
rlabel metal1 1 -826 1 -826 1 P3
rlabel metal1 1 -833 1 -833 1 G2
rlabel metal1 488 -752 488 -752 1 G3
<< end >>
