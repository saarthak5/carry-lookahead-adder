magic
tech scmos
timestamp 1732089451
<< nwell >>
rect 14 110 98 147
rect 14 27 38 64
rect 14 -40 98 -3
rect 14 -123 38 -86
rect 14 -190 98 -153
rect 14 -273 38 -236
rect 14 -340 98 -303
rect 14 -423 38 -386
<< ntransistor >>
rect 25 91 27 101
rect 25 8 27 18
rect 49 8 51 18
rect 66 8 68 18
rect 79 8 81 18
rect 96 8 98 18
rect 25 -59 27 -49
rect 25 -142 27 -132
rect 49 -142 51 -132
rect 66 -142 68 -132
rect 79 -142 81 -132
rect 96 -142 98 -132
rect 25 -209 27 -199
rect 25 -292 27 -282
rect 49 -292 51 -282
rect 66 -292 68 -282
rect 79 -292 81 -282
rect 96 -292 98 -282
rect 25 -359 27 -349
rect 25 -442 27 -432
rect 49 -442 51 -432
rect 66 -442 68 -432
rect 79 -442 81 -432
rect 96 -442 98 -432
<< ptransistor >>
rect 25 116 27 136
rect 49 116 51 136
rect 63 116 65 136
rect 71 116 73 136
rect 85 116 87 136
rect 25 33 27 53
rect 25 -34 27 -14
rect 49 -34 51 -14
rect 63 -34 65 -14
rect 71 -34 73 -14
rect 85 -34 87 -14
rect 25 -117 27 -97
rect 25 -184 27 -164
rect 49 -184 51 -164
rect 63 -184 65 -164
rect 71 -184 73 -164
rect 85 -184 87 -164
rect 25 -267 27 -247
rect 25 -334 27 -314
rect 49 -334 51 -314
rect 63 -334 65 -314
rect 71 -334 73 -314
rect 85 -334 87 -314
rect 25 -417 27 -397
<< ndiffusion >>
rect 24 91 25 101
rect 27 91 28 101
rect 24 8 25 18
rect 27 8 28 18
rect 48 8 49 18
rect 51 8 52 18
rect 65 8 66 18
rect 68 8 71 18
rect 75 8 79 18
rect 81 8 82 18
rect 95 8 96 18
rect 98 8 99 18
rect 24 -59 25 -49
rect 27 -59 28 -49
rect 24 -142 25 -132
rect 27 -142 28 -132
rect 48 -142 49 -132
rect 51 -142 52 -132
rect 65 -142 66 -132
rect 68 -142 71 -132
rect 75 -142 79 -132
rect 81 -142 82 -132
rect 95 -142 96 -132
rect 98 -142 99 -132
rect 24 -209 25 -199
rect 27 -209 28 -199
rect 24 -292 25 -282
rect 27 -292 28 -282
rect 48 -292 49 -282
rect 51 -292 52 -282
rect 65 -292 66 -282
rect 68 -292 71 -282
rect 75 -292 79 -282
rect 81 -292 82 -282
rect 95 -292 96 -282
rect 98 -292 99 -282
rect 24 -359 25 -349
rect 27 -359 28 -349
rect 24 -442 25 -432
rect 27 -442 28 -432
rect 48 -442 49 -432
rect 51 -442 52 -432
rect 65 -442 66 -432
rect 68 -442 71 -432
rect 75 -442 79 -432
rect 81 -442 82 -432
rect 95 -442 96 -432
rect 98 -442 99 -432
<< pdiffusion >>
rect 24 116 25 136
rect 27 116 28 136
rect 48 116 49 136
rect 51 116 63 136
rect 65 116 66 136
rect 70 116 71 136
rect 73 116 85 136
rect 87 116 88 136
rect 24 33 25 53
rect 27 33 28 53
rect 24 -34 25 -14
rect 27 -34 28 -14
rect 48 -34 49 -14
rect 51 -34 63 -14
rect 65 -34 66 -14
rect 70 -34 71 -14
rect 73 -34 85 -14
rect 87 -34 88 -14
rect 24 -117 25 -97
rect 27 -117 28 -97
rect 24 -184 25 -164
rect 27 -184 28 -164
rect 48 -184 49 -164
rect 51 -184 63 -164
rect 65 -184 66 -164
rect 70 -184 71 -164
rect 73 -184 85 -164
rect 87 -184 88 -164
rect 24 -267 25 -247
rect 27 -267 28 -247
rect 24 -334 25 -314
rect 27 -334 28 -314
rect 48 -334 49 -314
rect 51 -334 63 -314
rect 65 -334 66 -314
rect 70 -334 71 -314
rect 73 -334 85 -314
rect 87 -334 88 -314
rect 24 -417 25 -397
rect 27 -417 28 -397
<< ndcontact >>
rect 20 91 24 101
rect 28 91 32 101
rect 20 8 24 18
rect 28 8 32 18
rect 44 8 48 18
rect 52 8 56 18
rect 71 8 75 18
rect 82 8 86 18
rect 99 8 103 18
rect 20 -59 24 -49
rect 28 -59 32 -49
rect 20 -142 24 -132
rect 28 -142 32 -132
rect 44 -142 48 -132
rect 52 -142 56 -132
rect 71 -142 75 -132
rect 82 -142 86 -132
rect 99 -142 103 -132
rect 20 -209 24 -199
rect 28 -209 32 -199
rect 20 -292 24 -282
rect 28 -292 32 -282
rect 44 -292 48 -282
rect 52 -292 56 -282
rect 71 -292 75 -282
rect 82 -292 86 -282
rect 99 -292 103 -282
rect 20 -359 24 -349
rect 28 -359 32 -349
rect 20 -442 24 -432
rect 28 -442 32 -432
rect 44 -442 48 -432
rect 52 -442 56 -432
rect 71 -442 75 -432
rect 82 -442 86 -432
rect 99 -442 103 -432
<< pdcontact >>
rect 20 116 24 136
rect 28 116 32 136
rect 44 116 48 136
rect 66 116 70 136
rect 88 116 92 136
rect 20 33 24 53
rect 28 33 32 53
rect 20 -34 24 -14
rect 28 -34 32 -14
rect 44 -34 48 -14
rect 66 -34 70 -14
rect 88 -34 92 -14
rect 20 -117 24 -97
rect 28 -117 32 -97
rect 20 -184 24 -164
rect 28 -184 32 -164
rect 44 -184 48 -164
rect 66 -184 70 -164
rect 88 -184 92 -164
rect 20 -267 24 -247
rect 28 -267 32 -247
rect 20 -334 24 -314
rect 28 -334 32 -314
rect 44 -334 48 -314
rect 66 -334 70 -314
rect 88 -334 92 -314
rect 20 -417 24 -397
rect 28 -417 32 -397
<< psubstratepcontact >>
rect 24 0 28 4
rect 24 -150 28 -146
rect 24 -300 28 -296
rect 24 -450 28 -446
<< nsubstratencontact >>
rect 24 140 28 144
rect 24 57 28 61
rect 24 -10 28 -6
rect 24 -93 28 -89
rect 24 -160 28 -156
rect 24 -243 28 -239
rect 24 -310 28 -306
rect 24 -393 28 -389
<< polysilicon >>
rect 25 136 27 139
rect 49 136 51 139
rect 63 136 65 139
rect 71 136 73 139
rect 85 136 87 139
rect 25 101 27 116
rect 25 88 27 91
rect 25 53 27 56
rect 25 18 27 33
rect 49 18 51 116
rect 63 45 65 116
rect 58 43 65 45
rect 58 30 60 43
rect 58 28 65 30
rect 63 21 65 28
rect 71 21 73 116
rect 85 21 87 116
rect 63 19 68 21
rect 71 19 81 21
rect 85 19 98 21
rect 66 18 68 19
rect 79 18 81 19
rect 96 18 98 19
rect 25 5 27 8
rect 49 5 51 8
rect 66 5 68 8
rect 79 5 81 8
rect 96 5 98 8
rect 25 -14 27 -11
rect 49 -14 51 -11
rect 63 -14 65 -11
rect 71 -14 73 -11
rect 85 -14 87 -11
rect 25 -49 27 -34
rect 25 -62 27 -59
rect 25 -97 27 -94
rect 25 -132 27 -117
rect 49 -132 51 -34
rect 63 -105 65 -34
rect 58 -107 65 -105
rect 58 -120 60 -107
rect 58 -122 65 -120
rect 63 -129 65 -122
rect 71 -129 73 -34
rect 85 -129 87 -34
rect 63 -131 68 -129
rect 71 -131 81 -129
rect 85 -131 98 -129
rect 66 -132 68 -131
rect 79 -132 81 -131
rect 96 -132 98 -131
rect 25 -145 27 -142
rect 49 -145 51 -142
rect 66 -145 68 -142
rect 79 -145 81 -142
rect 96 -145 98 -142
rect 25 -164 27 -161
rect 49 -164 51 -161
rect 63 -164 65 -161
rect 71 -164 73 -161
rect 85 -164 87 -161
rect 25 -199 27 -184
rect 25 -212 27 -209
rect 25 -247 27 -244
rect 25 -282 27 -267
rect 49 -282 51 -184
rect 63 -255 65 -184
rect 58 -257 65 -255
rect 58 -270 60 -257
rect 58 -272 65 -270
rect 63 -279 65 -272
rect 71 -279 73 -184
rect 85 -279 87 -184
rect 63 -281 68 -279
rect 71 -281 81 -279
rect 85 -281 98 -279
rect 66 -282 68 -281
rect 79 -282 81 -281
rect 96 -282 98 -281
rect 25 -295 27 -292
rect 49 -295 51 -292
rect 66 -295 68 -292
rect 79 -295 81 -292
rect 96 -295 98 -292
rect 25 -314 27 -311
rect 49 -314 51 -311
rect 63 -314 65 -311
rect 71 -314 73 -311
rect 85 -314 87 -311
rect 25 -349 27 -334
rect 25 -362 27 -359
rect 25 -397 27 -394
rect 25 -432 27 -417
rect 49 -432 51 -334
rect 63 -405 65 -334
rect 58 -407 65 -405
rect 58 -420 60 -407
rect 58 -422 65 -420
rect 63 -429 65 -422
rect 71 -429 73 -334
rect 85 -429 87 -334
rect 63 -431 68 -429
rect 71 -431 81 -429
rect 85 -431 98 -429
rect 66 -432 68 -431
rect 79 -432 81 -431
rect 96 -432 98 -431
rect 25 -445 27 -442
rect 49 -445 51 -442
rect 66 -445 68 -442
rect 79 -445 81 -442
rect 96 -445 98 -442
<< polycontact >>
rect 21 105 25 109
rect 45 105 49 109
rect 21 22 25 26
rect 59 76 63 80
rect 21 -45 25 -41
rect 45 -45 49 -41
rect 21 -128 25 -124
rect 59 -74 63 -70
rect 21 -195 25 -191
rect 45 -195 49 -191
rect 21 -278 25 -274
rect 59 -224 63 -220
rect 21 -345 25 -341
rect 45 -345 49 -341
rect 21 -428 25 -424
rect 59 -374 63 -370
<< metal1 >>
rect 14 144 38 146
rect 14 140 24 144
rect 28 140 38 144
rect 43 140 92 146
rect 20 136 24 140
rect 44 136 48 140
rect 88 136 92 140
rect 28 109 32 116
rect 0 105 21 109
rect 28 105 45 109
rect 0 79 4 105
rect 28 101 32 105
rect 20 87 24 91
rect 12 82 24 87
rect 27 83 57 87
rect 27 79 31 83
rect 0 75 31 79
rect 34 76 59 80
rect 34 71 38 76
rect 66 73 70 116
rect 7 67 38 71
rect 44 69 103 73
rect 7 26 11 67
rect 14 61 33 63
rect 14 57 24 61
rect 28 57 33 61
rect 20 53 24 57
rect 28 26 32 33
rect 0 22 21 26
rect 28 21 33 26
rect 28 18 32 21
rect 44 18 48 69
rect 52 21 86 25
rect 52 18 56 21
rect 82 18 86 21
rect 99 18 103 69
rect 20 5 24 8
rect 12 0 24 5
rect 71 4 75 8
rect 28 0 75 4
rect 14 -6 38 -4
rect 14 -10 24 -6
rect 28 -10 38 -6
rect 43 -10 92 -4
rect 20 -14 24 -10
rect 44 -14 48 -10
rect 88 -14 92 -10
rect 28 -41 32 -34
rect 0 -45 21 -41
rect 28 -45 45 -41
rect 0 -71 4 -45
rect 28 -49 32 -45
rect 20 -63 24 -59
rect 12 -68 24 -63
rect 27 -67 57 -63
rect 27 -71 31 -67
rect 0 -75 31 -71
rect 34 -74 59 -70
rect 34 -79 38 -74
rect 66 -77 70 -34
rect 7 -83 38 -79
rect 44 -81 103 -77
rect 7 -124 11 -83
rect 14 -89 33 -87
rect 14 -93 24 -89
rect 28 -93 33 -89
rect 20 -97 24 -93
rect 28 -124 32 -117
rect 0 -128 21 -124
rect 28 -129 33 -124
rect 28 -132 32 -129
rect 44 -132 48 -81
rect 52 -129 86 -125
rect 52 -132 56 -129
rect 82 -132 86 -129
rect 99 -132 103 -81
rect 20 -145 24 -142
rect 12 -150 24 -145
rect 71 -146 75 -142
rect 28 -150 75 -146
rect 14 -156 38 -154
rect 14 -160 24 -156
rect 28 -160 38 -156
rect 43 -160 92 -154
rect 20 -164 24 -160
rect 44 -164 48 -160
rect 88 -164 92 -160
rect 28 -191 32 -184
rect 0 -195 21 -191
rect 28 -195 45 -191
rect 0 -221 4 -195
rect 28 -199 32 -195
rect 20 -213 24 -209
rect 12 -218 24 -213
rect 27 -217 57 -213
rect 27 -221 31 -217
rect 0 -225 31 -221
rect 34 -224 59 -220
rect 34 -229 38 -224
rect 66 -227 70 -184
rect 7 -233 38 -229
rect 44 -231 103 -227
rect 7 -274 11 -233
rect 14 -239 33 -237
rect 14 -243 24 -239
rect 28 -243 33 -239
rect 20 -247 24 -243
rect 28 -274 32 -267
rect 0 -278 21 -274
rect 28 -279 33 -274
rect 28 -282 32 -279
rect 44 -282 48 -231
rect 52 -279 86 -275
rect 52 -282 56 -279
rect 82 -282 86 -279
rect 99 -282 103 -231
rect 20 -295 24 -292
rect 12 -300 24 -295
rect 71 -296 75 -292
rect 28 -300 75 -296
rect 14 -306 38 -304
rect 14 -310 24 -306
rect 28 -310 38 -306
rect 43 -310 92 -304
rect 20 -314 24 -310
rect 44 -314 48 -310
rect 88 -314 92 -310
rect 28 -341 32 -334
rect 0 -345 21 -341
rect 28 -345 45 -341
rect 0 -371 4 -345
rect 28 -349 32 -345
rect 20 -363 24 -359
rect 12 -368 24 -363
rect 27 -367 57 -363
rect 27 -371 31 -367
rect 0 -375 31 -371
rect 34 -374 59 -370
rect 34 -379 38 -374
rect 66 -377 70 -334
rect 7 -383 38 -379
rect 44 -381 103 -377
rect 7 -424 11 -383
rect 14 -389 33 -387
rect 14 -393 24 -389
rect 28 -393 33 -389
rect 20 -397 24 -393
rect 28 -424 32 -417
rect 0 -428 21 -424
rect 28 -429 33 -424
rect 28 -432 32 -429
rect 44 -432 48 -381
rect 52 -429 86 -425
rect 52 -432 56 -429
rect 82 -432 86 -429
rect 99 -432 103 -381
rect 20 -445 24 -442
rect 12 -450 24 -445
rect 71 -446 75 -442
rect 28 -450 75 -446
<< m2contact >>
rect 38 140 43 146
rect 7 82 12 87
rect 57 83 62 88
rect 33 57 38 63
rect 33 21 38 26
rect 7 0 12 5
rect 38 -10 43 -4
rect 7 -68 12 -63
rect 57 -67 62 -62
rect 33 -93 38 -87
rect 33 -129 38 -124
rect 7 -150 12 -145
rect 38 -160 43 -154
rect 7 -218 12 -213
rect 57 -217 62 -212
rect 33 -243 38 -237
rect 33 -279 38 -274
rect 7 -300 12 -295
rect 38 -310 43 -304
rect 7 -368 12 -363
rect 57 -367 62 -362
rect 33 -393 38 -387
rect 33 -429 38 -424
rect 7 -450 12 -445
<< pm12contact >>
rect 80 83 85 88
rect 66 34 71 39
rect 80 -67 85 -62
rect 66 -116 71 -111
rect 80 -217 85 -212
rect 66 -266 71 -261
rect 80 -367 85 -362
rect 66 -416 71 -411
<< ndm12contact >>
rect 60 8 65 18
rect 90 8 95 18
rect 60 -142 65 -132
rect 90 -142 95 -132
rect 60 -292 65 -282
rect 90 -292 95 -282
rect 60 -442 65 -432
rect 90 -442 95 -432
<< metal2 >>
rect 7 5 12 82
rect 38 57 43 140
rect 62 83 80 88
rect 38 34 66 39
rect 38 21 43 34
rect 60 21 95 25
rect 60 18 65 21
rect 90 18 95 21
rect 7 -145 12 -68
rect 38 -93 43 -10
rect 62 -67 80 -62
rect 38 -116 66 -111
rect 38 -129 43 -116
rect 60 -129 95 -125
rect 60 -132 65 -129
rect 90 -132 95 -129
rect 7 -295 12 -218
rect 38 -243 43 -160
rect 62 -217 80 -212
rect 38 -266 66 -261
rect 38 -279 43 -266
rect 60 -279 95 -275
rect 60 -282 65 -279
rect 90 -282 95 -279
rect 7 -445 12 -368
rect 38 -393 43 -310
rect 62 -367 80 -362
rect 38 -416 66 -411
rect 38 -429 43 -416
rect 60 -429 95 -425
rect 60 -432 65 -429
rect 90 -432 95 -429
<< labels >>
rlabel metal1 17 143 17 143 4 vdd
rlabel metal1 16 2 16 2 2 gnd
rlabel metal1 101 71 101 71 7 S0
rlabel metal1 15 107 15 107 1 P0
rlabel metal1 15 24 15 24 1 Cin
rlabel metal1 17 -7 17 -7 4 vdd
rlabel metal1 16 -148 16 -148 2 gnd
rlabel metal1 17 -157 17 -157 4 vdd
rlabel metal1 16 -298 16 -298 2 gnd
rlabel metal1 17 -307 17 -307 4 vdd
rlabel metal1 16 -448 16 -448 2 gnd
rlabel metal1 15 -43 15 -43 1 P1
rlabel metal1 15 -126 15 -126 1 C1
rlabel metal1 15 -193 15 -193 1 P2
rlabel metal1 15 -276 15 -276 1 C2
rlabel metal1 15 -343 15 -343 1 P3
rlabel metal1 15 -426 15 -426 1 C3
rlabel metal1 101 -379 101 -379 7 S3
rlabel metal1 101 -229 101 -229 7 S2
rlabel metal1 101 -79 101 -79 7 S1
<< end >>
