magic
tech scmos
timestamp 1732080839
<< nwell >>
rect 14 110 98 147
rect 14 27 38 64
rect 4 -40 66 -3
rect 14 -114 98 -77
rect 14 -197 38 -160
rect 4 -264 66 -227
rect 14 -338 98 -301
rect 14 -421 38 -384
rect 4 -488 66 -451
rect 14 -562 98 -525
rect 14 -645 38 -608
rect 4 -712 66 -675
<< ntransistor >>
rect 25 91 27 101
rect 25 8 27 18
rect 49 8 51 18
rect 66 8 68 18
rect 79 8 81 18
rect 96 8 98 18
rect 15 -66 17 -56
rect 29 -66 31 -56
rect 53 -66 55 -56
rect 25 -133 27 -123
rect 25 -216 27 -206
rect 49 -216 51 -206
rect 66 -216 68 -206
rect 79 -216 81 -206
rect 96 -216 98 -206
rect 15 -290 17 -280
rect 29 -290 31 -280
rect 53 -290 55 -280
rect 25 -357 27 -347
rect 25 -440 27 -430
rect 49 -440 51 -430
rect 66 -440 68 -430
rect 79 -440 81 -430
rect 96 -440 98 -430
rect 15 -514 17 -504
rect 29 -514 31 -504
rect 53 -514 55 -504
rect 25 -581 27 -571
rect 25 -664 27 -654
rect 49 -664 51 -654
rect 66 -664 68 -654
rect 79 -664 81 -654
rect 96 -664 98 -654
rect 15 -738 17 -728
rect 29 -738 31 -728
rect 53 -738 55 -728
<< ptransistor >>
rect 25 116 27 136
rect 49 116 51 136
rect 63 116 65 136
rect 71 116 73 136
rect 85 116 87 136
rect 25 33 27 53
rect 15 -34 17 -14
rect 29 -34 31 -14
rect 53 -34 55 -14
rect 25 -108 27 -88
rect 49 -108 51 -88
rect 63 -108 65 -88
rect 71 -108 73 -88
rect 85 -108 87 -88
rect 25 -191 27 -171
rect 15 -258 17 -238
rect 29 -258 31 -238
rect 53 -258 55 -238
rect 25 -332 27 -312
rect 49 -332 51 -312
rect 63 -332 65 -312
rect 71 -332 73 -312
rect 85 -332 87 -312
rect 25 -415 27 -395
rect 15 -482 17 -462
rect 29 -482 31 -462
rect 53 -482 55 -462
rect 25 -556 27 -536
rect 49 -556 51 -536
rect 63 -556 65 -536
rect 71 -556 73 -536
rect 85 -556 87 -536
rect 25 -639 27 -619
rect 15 -706 17 -686
rect 29 -706 31 -686
rect 53 -706 55 -686
<< ndiffusion >>
rect 24 91 25 101
rect 27 91 28 101
rect 24 8 25 18
rect 27 8 28 18
rect 48 8 49 18
rect 51 8 52 18
rect 65 8 66 18
rect 68 8 71 18
rect 75 8 79 18
rect 81 8 82 18
rect 95 8 96 18
rect 98 8 99 18
rect 14 -66 15 -56
rect 17 -66 29 -56
rect 31 -66 32 -56
rect 52 -66 53 -56
rect 55 -66 56 -56
rect 24 -133 25 -123
rect 27 -133 28 -123
rect 24 -216 25 -206
rect 27 -216 28 -206
rect 48 -216 49 -206
rect 51 -216 52 -206
rect 65 -216 66 -206
rect 68 -216 71 -206
rect 75 -216 79 -206
rect 81 -216 82 -206
rect 95 -216 96 -206
rect 98 -216 99 -206
rect 14 -290 15 -280
rect 17 -290 29 -280
rect 31 -290 32 -280
rect 52 -290 53 -280
rect 55 -290 56 -280
rect 24 -357 25 -347
rect 27 -357 28 -347
rect 24 -440 25 -430
rect 27 -440 28 -430
rect 48 -440 49 -430
rect 51 -440 52 -430
rect 65 -440 66 -430
rect 68 -440 71 -430
rect 75 -440 79 -430
rect 81 -440 82 -430
rect 95 -440 96 -430
rect 98 -440 99 -430
rect 14 -514 15 -504
rect 17 -514 29 -504
rect 31 -514 32 -504
rect 52 -514 53 -504
rect 55 -514 56 -504
rect 24 -581 25 -571
rect 27 -581 28 -571
rect 24 -664 25 -654
rect 27 -664 28 -654
rect 48 -664 49 -654
rect 51 -664 52 -654
rect 65 -664 66 -654
rect 68 -664 71 -654
rect 75 -664 79 -654
rect 81 -664 82 -654
rect 95 -664 96 -654
rect 98 -664 99 -654
rect 14 -738 15 -728
rect 17 -738 29 -728
rect 31 -738 32 -728
rect 52 -738 53 -728
rect 55 -738 56 -728
<< pdiffusion >>
rect 24 116 25 136
rect 27 116 28 136
rect 48 116 49 136
rect 51 116 63 136
rect 65 116 66 136
rect 70 116 71 136
rect 73 116 85 136
rect 87 116 88 136
rect 24 33 25 53
rect 27 33 28 53
rect 14 -34 15 -14
rect 17 -34 21 -14
rect 25 -34 29 -14
rect 31 -34 32 -14
rect 52 -34 53 -14
rect 55 -34 56 -14
rect 24 -108 25 -88
rect 27 -108 28 -88
rect 48 -108 49 -88
rect 51 -108 63 -88
rect 65 -108 66 -88
rect 70 -108 71 -88
rect 73 -108 85 -88
rect 87 -108 88 -88
rect 24 -191 25 -171
rect 27 -191 28 -171
rect 14 -258 15 -238
rect 17 -258 21 -238
rect 25 -258 29 -238
rect 31 -258 32 -238
rect 52 -258 53 -238
rect 55 -258 56 -238
rect 24 -332 25 -312
rect 27 -332 28 -312
rect 48 -332 49 -312
rect 51 -332 63 -312
rect 65 -332 66 -312
rect 70 -332 71 -312
rect 73 -332 85 -312
rect 87 -332 88 -312
rect 24 -415 25 -395
rect 27 -415 28 -395
rect 14 -482 15 -462
rect 17 -482 21 -462
rect 25 -482 29 -462
rect 31 -482 32 -462
rect 52 -482 53 -462
rect 55 -482 56 -462
rect 24 -556 25 -536
rect 27 -556 28 -536
rect 48 -556 49 -536
rect 51 -556 63 -536
rect 65 -556 66 -536
rect 70 -556 71 -536
rect 73 -556 85 -536
rect 87 -556 88 -536
rect 24 -639 25 -619
rect 27 -639 28 -619
rect 14 -706 15 -686
rect 17 -706 21 -686
rect 25 -706 29 -686
rect 31 -706 32 -686
rect 52 -706 53 -686
rect 55 -706 56 -686
<< ndcontact >>
rect 20 91 24 101
rect 28 91 32 101
rect 20 8 24 18
rect 28 8 32 18
rect 44 8 48 18
rect 52 8 56 18
rect 71 8 75 18
rect 82 8 86 18
rect 99 8 103 18
rect 10 -66 14 -56
rect 32 -66 36 -56
rect 48 -66 52 -56
rect 56 -66 60 -56
rect 20 -133 24 -123
rect 28 -133 32 -123
rect 20 -216 24 -206
rect 28 -216 32 -206
rect 44 -216 48 -206
rect 52 -216 56 -206
rect 71 -216 75 -206
rect 82 -216 86 -206
rect 99 -216 103 -206
rect 10 -290 14 -280
rect 32 -290 36 -280
rect 48 -290 52 -280
rect 56 -290 60 -280
rect 20 -357 24 -347
rect 28 -357 32 -347
rect 20 -440 24 -430
rect 28 -440 32 -430
rect 44 -440 48 -430
rect 52 -440 56 -430
rect 71 -440 75 -430
rect 82 -440 86 -430
rect 99 -440 103 -430
rect 10 -514 14 -504
rect 32 -514 36 -504
rect 48 -514 52 -504
rect 56 -514 60 -504
rect 20 -581 24 -571
rect 28 -581 32 -571
rect 20 -664 24 -654
rect 28 -664 32 -654
rect 44 -664 48 -654
rect 52 -664 56 -654
rect 71 -664 75 -654
rect 82 -664 86 -654
rect 99 -664 103 -654
rect 10 -738 14 -728
rect 32 -738 36 -728
rect 48 -738 52 -728
rect 56 -738 60 -728
<< pdcontact >>
rect 20 116 24 136
rect 28 116 32 136
rect 44 116 48 136
rect 66 116 70 136
rect 88 116 92 136
rect 20 33 24 53
rect 28 33 32 53
rect 10 -34 14 -14
rect 21 -34 25 -14
rect 32 -34 36 -14
rect 48 -34 52 -14
rect 56 -34 60 -14
rect 20 -108 24 -88
rect 28 -108 32 -88
rect 44 -108 48 -88
rect 66 -108 70 -88
rect 88 -108 92 -88
rect 20 -191 24 -171
rect 28 -191 32 -171
rect 10 -258 14 -238
rect 21 -258 25 -238
rect 32 -258 36 -238
rect 48 -258 52 -238
rect 56 -258 60 -238
rect 20 -332 24 -312
rect 28 -332 32 -312
rect 44 -332 48 -312
rect 66 -332 70 -312
rect 88 -332 92 -312
rect 20 -415 24 -395
rect 28 -415 32 -395
rect 10 -482 14 -462
rect 21 -482 25 -462
rect 32 -482 36 -462
rect 48 -482 52 -462
rect 56 -482 60 -462
rect 20 -556 24 -536
rect 28 -556 32 -536
rect 44 -556 48 -536
rect 66 -556 70 -536
rect 88 -556 92 -536
rect 20 -639 24 -619
rect 28 -639 32 -619
rect 10 -706 14 -686
rect 21 -706 25 -686
rect 32 -706 36 -686
rect 48 -706 52 -686
rect 56 -706 60 -686
<< psubstratepcontact >>
rect 24 0 28 4
rect 52 -74 56 -70
rect 24 -224 28 -220
rect 52 -298 56 -294
rect 24 -448 28 -444
rect 52 -522 56 -518
rect 24 -672 28 -668
rect 52 -746 56 -742
<< nsubstratencontact >>
rect 24 140 28 144
rect 24 57 28 61
rect 52 -10 56 -6
rect 24 -84 28 -80
rect 24 -167 28 -163
rect 52 -234 56 -230
rect 24 -308 28 -304
rect 24 -391 28 -387
rect 52 -458 56 -454
rect 24 -532 28 -528
rect 24 -615 28 -611
rect 52 -682 56 -678
<< polysilicon >>
rect 25 136 27 139
rect 49 136 51 139
rect 63 136 65 139
rect 71 136 73 139
rect 85 136 87 139
rect 25 101 27 116
rect 25 88 27 91
rect 25 53 27 56
rect 25 18 27 33
rect 49 18 51 116
rect 63 45 65 116
rect 58 43 65 45
rect 58 30 60 43
rect 58 28 65 30
rect 63 21 65 28
rect 71 21 73 116
rect 85 21 87 116
rect 63 19 68 21
rect 71 19 81 21
rect 85 19 98 21
rect 66 18 68 19
rect 79 18 81 19
rect 96 18 98 19
rect 25 5 27 8
rect 49 5 51 8
rect 66 5 68 8
rect 79 5 81 8
rect 96 5 98 8
rect 15 -14 17 -11
rect 29 -14 31 -11
rect 53 -14 55 -11
rect 15 -56 17 -34
rect 29 -56 31 -34
rect 53 -56 55 -34
rect 15 -69 17 -66
rect 29 -69 31 -66
rect 53 -69 55 -66
rect 25 -88 27 -85
rect 49 -88 51 -85
rect 63 -88 65 -85
rect 71 -88 73 -85
rect 85 -88 87 -85
rect 25 -123 27 -108
rect 25 -136 27 -133
rect 25 -171 27 -168
rect 25 -206 27 -191
rect 49 -206 51 -108
rect 63 -179 65 -108
rect 58 -181 65 -179
rect 58 -194 60 -181
rect 58 -196 65 -194
rect 63 -203 65 -196
rect 71 -203 73 -108
rect 85 -203 87 -108
rect 63 -205 68 -203
rect 71 -205 81 -203
rect 85 -205 98 -203
rect 66 -206 68 -205
rect 79 -206 81 -205
rect 96 -206 98 -205
rect 25 -219 27 -216
rect 49 -219 51 -216
rect 66 -219 68 -216
rect 79 -219 81 -216
rect 96 -219 98 -216
rect 15 -238 17 -235
rect 29 -238 31 -235
rect 53 -238 55 -235
rect 15 -280 17 -258
rect 29 -280 31 -258
rect 53 -280 55 -258
rect 15 -293 17 -290
rect 29 -293 31 -290
rect 53 -293 55 -290
rect 25 -312 27 -309
rect 49 -312 51 -309
rect 63 -312 65 -309
rect 71 -312 73 -309
rect 85 -312 87 -309
rect 25 -347 27 -332
rect 25 -360 27 -357
rect 25 -395 27 -392
rect 25 -430 27 -415
rect 49 -430 51 -332
rect 63 -403 65 -332
rect 58 -405 65 -403
rect 58 -418 60 -405
rect 58 -420 65 -418
rect 63 -427 65 -420
rect 71 -427 73 -332
rect 85 -427 87 -332
rect 63 -429 68 -427
rect 71 -429 81 -427
rect 85 -429 98 -427
rect 66 -430 68 -429
rect 79 -430 81 -429
rect 96 -430 98 -429
rect 25 -443 27 -440
rect 49 -443 51 -440
rect 66 -443 68 -440
rect 79 -443 81 -440
rect 96 -443 98 -440
rect 15 -462 17 -459
rect 29 -462 31 -459
rect 53 -462 55 -459
rect 15 -504 17 -482
rect 29 -504 31 -482
rect 53 -504 55 -482
rect 15 -517 17 -514
rect 29 -517 31 -514
rect 53 -517 55 -514
rect 25 -536 27 -533
rect 49 -536 51 -533
rect 63 -536 65 -533
rect 71 -536 73 -533
rect 85 -536 87 -533
rect 25 -571 27 -556
rect 25 -584 27 -581
rect 25 -619 27 -616
rect 25 -654 27 -639
rect 49 -654 51 -556
rect 63 -627 65 -556
rect 58 -629 65 -627
rect 58 -642 60 -629
rect 58 -644 65 -642
rect 63 -651 65 -644
rect 71 -651 73 -556
rect 85 -651 87 -556
rect 63 -653 68 -651
rect 71 -653 81 -651
rect 85 -653 98 -651
rect 66 -654 68 -653
rect 79 -654 81 -653
rect 96 -654 98 -653
rect 25 -667 27 -664
rect 49 -667 51 -664
rect 66 -667 68 -664
rect 79 -667 81 -664
rect 96 -667 98 -664
rect 15 -686 17 -683
rect 29 -686 31 -683
rect 53 -686 55 -683
rect 15 -728 17 -706
rect 29 -728 31 -706
rect 53 -728 55 -706
rect 15 -741 17 -738
rect 29 -741 31 -738
rect 53 -741 55 -738
<< polycontact >>
rect 21 105 25 109
rect 45 105 49 109
rect 21 22 25 26
rect 59 76 63 80
rect 11 -45 15 -41
rect 25 -52 29 -48
rect 49 -45 53 -41
rect 21 -119 25 -115
rect 45 -119 49 -115
rect 21 -202 25 -198
rect 59 -148 63 -144
rect 11 -269 15 -265
rect 25 -276 29 -272
rect 49 -269 53 -265
rect 21 -343 25 -339
rect 45 -343 49 -339
rect 21 -426 25 -422
rect 59 -372 63 -368
rect 11 -493 15 -489
rect 25 -500 29 -496
rect 49 -493 53 -489
rect 21 -567 25 -563
rect 45 -567 49 -563
rect 21 -650 25 -646
rect 59 -596 63 -592
rect 11 -717 15 -713
rect 25 -724 29 -720
rect 49 -717 53 -713
<< metal1 >>
rect 14 144 38 146
rect 14 140 24 144
rect 28 140 38 144
rect 43 140 87 146
rect 20 136 24 140
rect 44 136 48 140
rect 88 136 92 140
rect 28 109 32 116
rect 0 105 21 109
rect 28 105 45 109
rect 0 79 4 105
rect 28 101 32 105
rect 20 87 24 91
rect 12 82 24 87
rect 27 83 57 87
rect 27 79 31 83
rect -24 75 31 79
rect 34 76 59 80
rect -24 74 -5 75
rect -24 22 -19 27
rect -9 -48 -5 74
rect 34 71 38 76
rect 66 73 70 116
rect 7 67 38 71
rect 44 69 112 73
rect 7 26 11 67
rect 14 61 33 63
rect 14 57 24 61
rect 28 57 33 61
rect 20 53 24 57
rect 28 26 32 33
rect 3 22 21 26
rect 0 -41 4 22
rect 28 21 33 26
rect 28 18 32 21
rect 44 18 48 69
rect 52 21 86 25
rect 52 18 56 21
rect 82 18 86 21
rect 99 18 103 69
rect 20 5 24 8
rect 12 0 24 5
rect 71 4 75 8
rect 28 0 75 4
rect 10 -6 61 -4
rect 10 -10 52 -6
rect 56 -10 61 -6
rect 10 -14 14 -10
rect 32 -14 36 -10
rect 48 -14 52 -10
rect 21 -41 25 -34
rect 56 -41 60 -34
rect 0 -45 11 -41
rect 21 -45 49 -41
rect 56 -45 112 -41
rect -9 -52 25 -48
rect 32 -56 36 -45
rect 56 -56 60 -45
rect 10 -69 14 -66
rect 12 -70 14 -69
rect 48 -70 52 -66
rect 12 -74 52 -70
rect 14 -80 38 -78
rect 14 -84 24 -80
rect 28 -84 38 -80
rect 43 -84 87 -78
rect 20 -88 24 -84
rect 44 -88 48 -84
rect 88 -88 92 -84
rect 28 -115 32 -108
rect 0 -119 21 -115
rect 28 -119 45 -115
rect 0 -145 4 -119
rect 28 -123 32 -119
rect 20 -137 24 -133
rect 12 -142 24 -137
rect 27 -141 57 -137
rect 27 -145 31 -141
rect -24 -149 31 -145
rect 34 -148 59 -144
rect -24 -150 -5 -149
rect -24 -202 -19 -197
rect -9 -272 -5 -150
rect 34 -153 38 -148
rect 66 -151 70 -108
rect 7 -157 38 -153
rect 44 -155 112 -151
rect 7 -198 11 -157
rect 14 -163 33 -161
rect 14 -167 24 -163
rect 28 -167 33 -163
rect 20 -171 24 -167
rect 28 -198 32 -191
rect 3 -202 21 -198
rect 0 -265 4 -202
rect 28 -203 33 -198
rect 28 -206 32 -203
rect 44 -206 48 -155
rect 52 -203 86 -199
rect 52 -206 56 -203
rect 82 -206 86 -203
rect 99 -206 103 -155
rect 20 -219 24 -216
rect 12 -224 24 -219
rect 71 -220 75 -216
rect 28 -224 75 -220
rect 10 -230 61 -228
rect 10 -234 52 -230
rect 56 -234 61 -230
rect 10 -238 14 -234
rect 32 -238 36 -234
rect 48 -238 52 -234
rect 21 -265 25 -258
rect 56 -265 60 -258
rect 0 -269 11 -265
rect 21 -269 49 -265
rect 56 -269 112 -265
rect -9 -276 25 -272
rect 32 -280 36 -269
rect 56 -280 60 -269
rect 10 -293 14 -290
rect 12 -294 14 -293
rect 48 -294 52 -290
rect 12 -298 52 -294
rect 14 -304 38 -302
rect 14 -308 24 -304
rect 28 -308 38 -304
rect 43 -308 87 -302
rect 20 -312 24 -308
rect 44 -312 48 -308
rect 88 -312 92 -308
rect 28 -339 32 -332
rect 0 -343 21 -339
rect 28 -343 45 -339
rect 0 -369 4 -343
rect 28 -347 32 -343
rect 20 -361 24 -357
rect 12 -366 24 -361
rect 27 -365 57 -361
rect 27 -369 31 -365
rect -24 -373 31 -369
rect 34 -372 59 -368
rect -24 -374 -5 -373
rect -24 -426 -19 -421
rect -9 -496 -5 -374
rect 34 -377 38 -372
rect 66 -375 70 -332
rect 7 -381 38 -377
rect 44 -379 112 -375
rect 7 -422 11 -381
rect 14 -387 33 -385
rect 14 -391 24 -387
rect 28 -391 33 -387
rect 20 -395 24 -391
rect 28 -422 32 -415
rect 3 -426 21 -422
rect 0 -489 4 -426
rect 28 -427 33 -422
rect 28 -430 32 -427
rect 44 -430 48 -379
rect 52 -427 86 -423
rect 52 -430 56 -427
rect 82 -430 86 -427
rect 99 -430 103 -379
rect 20 -443 24 -440
rect 12 -448 24 -443
rect 71 -444 75 -440
rect 28 -448 75 -444
rect 10 -454 61 -452
rect 10 -458 52 -454
rect 56 -458 61 -454
rect 10 -462 14 -458
rect 32 -462 36 -458
rect 48 -462 52 -458
rect 21 -489 25 -482
rect 56 -489 60 -482
rect 0 -493 11 -489
rect 21 -493 49 -489
rect 56 -493 112 -489
rect -9 -500 25 -496
rect 32 -504 36 -493
rect 56 -504 60 -493
rect 10 -517 14 -514
rect 12 -518 14 -517
rect 48 -518 52 -514
rect 12 -522 52 -518
rect 14 -528 38 -526
rect 14 -532 24 -528
rect 28 -532 38 -528
rect 43 -532 87 -526
rect 20 -536 24 -532
rect 44 -536 48 -532
rect 88 -536 92 -532
rect 28 -563 32 -556
rect 0 -567 21 -563
rect 28 -567 45 -563
rect 0 -593 4 -567
rect 28 -571 32 -567
rect 20 -585 24 -581
rect 12 -590 24 -585
rect 27 -589 57 -585
rect 27 -593 31 -589
rect -24 -597 31 -593
rect 34 -596 59 -592
rect -24 -598 -5 -597
rect -24 -650 -19 -645
rect -9 -720 -5 -598
rect 34 -601 38 -596
rect 66 -599 70 -556
rect 7 -605 38 -601
rect 44 -603 112 -599
rect 7 -646 11 -605
rect 14 -611 33 -609
rect 14 -615 24 -611
rect 28 -615 33 -611
rect 20 -619 24 -615
rect 28 -646 32 -639
rect 3 -650 21 -646
rect 0 -713 4 -650
rect 28 -651 33 -646
rect 28 -654 32 -651
rect 44 -654 48 -603
rect 52 -651 86 -647
rect 52 -654 56 -651
rect 82 -654 86 -651
rect 99 -654 103 -603
rect 20 -667 24 -664
rect 12 -672 24 -667
rect 71 -668 75 -664
rect 28 -672 75 -668
rect 10 -678 61 -676
rect 10 -682 52 -678
rect 56 -682 61 -678
rect 10 -686 14 -682
rect 32 -686 36 -682
rect 48 -686 52 -682
rect 21 -713 25 -706
rect 56 -713 60 -706
rect 0 -717 11 -713
rect 21 -717 49 -713
rect 56 -717 112 -713
rect -9 -724 25 -720
rect 32 -728 36 -717
rect 56 -728 60 -717
rect 10 -741 14 -738
rect 12 -742 14 -741
rect 48 -742 52 -738
rect 12 -746 52 -742
<< m2contact >>
rect 38 140 43 146
rect 87 140 92 146
rect 7 82 12 87
rect 57 83 62 88
rect -19 22 -14 27
rect -2 22 3 27
rect 33 57 38 63
rect 33 21 38 26
rect 7 0 12 5
rect 61 -10 66 -4
rect 7 -74 12 -69
rect 38 -84 43 -78
rect 87 -84 92 -78
rect 7 -142 12 -137
rect 57 -141 62 -136
rect -19 -202 -14 -197
rect -2 -202 3 -197
rect 33 -167 38 -161
rect 33 -203 38 -198
rect 7 -224 12 -219
rect 61 -234 66 -228
rect 7 -298 12 -293
rect 38 -308 43 -302
rect 87 -308 92 -302
rect 7 -366 12 -361
rect 57 -365 62 -360
rect -19 -426 -14 -421
rect -2 -426 3 -421
rect 33 -391 38 -385
rect 33 -427 38 -422
rect 7 -448 12 -443
rect 61 -458 66 -452
rect 7 -522 12 -517
rect 38 -532 43 -526
rect 87 -532 92 -526
rect 7 -590 12 -585
rect 57 -589 62 -584
rect -19 -650 -14 -645
rect -2 -650 3 -645
rect 33 -615 38 -609
rect 33 -651 38 -646
rect 7 -672 12 -667
rect 61 -682 66 -676
rect 7 -746 12 -741
<< pm12contact >>
rect 80 83 85 88
rect 66 34 71 39
rect 80 -141 85 -136
rect 66 -190 71 -185
rect 80 -365 85 -360
rect 66 -414 71 -409
rect 80 -589 85 -584
rect 66 -638 71 -633
<< ndm12contact >>
rect 60 8 65 18
rect 90 8 95 18
rect 60 -216 65 -206
rect 90 -216 95 -206
rect 60 -440 65 -430
rect 90 -440 95 -430
rect 60 -664 65 -654
rect 90 -664 95 -654
<< metal2 >>
rect 92 140 108 146
rect -14 22 -2 27
rect 7 5 12 82
rect 38 57 43 140
rect 62 83 80 88
rect 38 34 66 39
rect 38 21 43 34
rect 60 21 95 25
rect 60 18 65 21
rect 90 18 95 21
rect 7 -69 12 0
rect 102 -4 108 140
rect 66 -10 108 -4
rect 7 -137 12 -74
rect 102 -78 108 -10
rect -14 -202 -2 -197
rect 7 -219 12 -142
rect 92 -84 108 -78
rect 38 -167 43 -84
rect 62 -141 80 -136
rect 38 -190 66 -185
rect 38 -203 43 -190
rect 60 -203 95 -199
rect 60 -206 65 -203
rect 90 -206 95 -203
rect 7 -293 12 -224
rect 102 -228 108 -84
rect 66 -234 108 -228
rect 7 -361 12 -298
rect 102 -302 108 -234
rect -14 -426 -2 -421
rect 7 -443 12 -366
rect 92 -308 108 -302
rect 38 -391 43 -308
rect 62 -365 80 -360
rect 38 -414 66 -409
rect 38 -427 43 -414
rect 60 -427 95 -423
rect 60 -430 65 -427
rect 90 -430 95 -427
rect 7 -517 12 -448
rect 102 -452 108 -308
rect 66 -458 108 -452
rect 7 -585 12 -522
rect 102 -526 108 -458
rect -14 -650 -2 -645
rect 7 -667 12 -590
rect 92 -532 108 -526
rect 38 -615 43 -532
rect 62 -589 80 -584
rect 38 -638 66 -633
rect 38 -651 43 -638
rect 60 -651 95 -647
rect 60 -654 65 -651
rect 90 -654 95 -651
rect 7 -741 12 -672
rect 102 -676 108 -532
rect 66 -682 108 -676
<< labels >>
rlabel metal1 16 143 16 143 5 vdd
rlabel metal1 -22 76 -22 76 3 A0
rlabel metal1 -23 24 -23 24 3 B0
rlabel metal1 111 71 111 71 7 P0
rlabel metal1 111 -43 111 -43 7 G0
rlabel metal1 -22 -148 -22 -148 3 A1
rlabel metal1 -22 -200 -22 -200 3 B1
rlabel metal1 111 -153 111 -153 7 P1
rlabel metal1 111 -267 111 -267 7 G1
rlabel metal1 -22 -372 -22 -372 3 A2
rlabel metal1 -23 -424 -23 -424 3 B2
rlabel metal1 111 -377 111 -377 7 P2
rlabel metal1 111 -491 111 -491 7 G2
rlabel metal1 -22 -596 -22 -596 3 A3
rlabel metal1 -23 -648 -23 -648 3 B3
rlabel metal1 111 -601 111 -601 7 P3
rlabel metal1 110 -715 110 -715 7 G3
rlabel metal1 35 -744 35 -744 1 gnd
<< end >>
