* SPICE3 file created from not.ext - technology: scmos

.include TSMC_180nm.txt
.param supply=1.8
.global gnd vdd
.option scale=0.09u

* source		nodes			value
*******************************************************************
vdd				vdd	gnd			'supply'
vin				in	gnd			pulse 0 'supply' 0 10p 10p 5n 10n

M1000 out in vdd vdd CMOSP w=20 l=2
+  ad=100 pd=50 as=100 ps=50
M1001 out in gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=50 ps=30
C0 in out 0.05fF
C1 vdd in 0.09fF
C2 gnd in 0.04fF
C3 vdd out 0.29fF
C4 gnd out 0.14fF
C5 gnd Gnd 0.08fF
C6 out Gnd 0.06fF
C7 in Gnd 0.14fF
C8 vdd Gnd 0.90fF

.control
tran 100p 20n
run

set hcopypscolor=1
set color0=white
set color1=black

set curplottitle='Saarthak-Sabharwal-2023102055-not-post'
plot V(out) V(in)+2
*hardcopy not.eps V(out) V(in)+2
.endc

.end
